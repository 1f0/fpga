`timescale 1ns / 1ps
module font_table (a,d);
    input  [12:0] a; // 8*8*128=2^3*2^3*2^7
    output        d; // font dot
    wire          rom [0:8191];
    assign        d = rom[a];

    assign rom[13'h0000] = 0;
    assign rom[13'h0001] = 0;
    assign rom[13'h0002] = 0;
    assign rom[13'h0003] = 0;
    assign rom[13'h0004] = 0;
    assign rom[13'h0005] = 0;
    assign rom[13'h0006] = 0;
    assign rom[13'h0007] = 0;
    assign rom[13'h0008] = 0;
    assign rom[13'h0009] = 0;
    assign rom[13'h000a] = 0;
    assign rom[13'h000b] = 0;
    assign rom[13'h000c] = 0;
    assign rom[13'h000d] = 0;
    assign rom[13'h000e] = 0;
    assign rom[13'h000f] = 0;
    assign rom[13'h0010] = 0;
    assign rom[13'h0011] = 0;
    assign rom[13'h0012] = 0;
    assign rom[13'h0013] = 0;
    assign rom[13'h0014] = 0;
    assign rom[13'h0015] = 0;
    assign rom[13'h0016] = 0;
    assign rom[13'h0017] = 0;
    assign rom[13'h0018] = 0;
    assign rom[13'h0019] = 0;
    assign rom[13'h001a] = 0;
    assign rom[13'h001b] = 0;
    assign rom[13'h001c] = 0;
    assign rom[13'h001d] = 0;
    assign rom[13'h001e] = 0;
    assign rom[13'h001f] = 0;
    assign rom[13'h0020] = 0;
    assign rom[13'h0021] = 0;
    assign rom[13'h0022] = 0;
    assign rom[13'h0023] = 0;
    assign rom[13'h0024] = 0;
    assign rom[13'h0025] = 0;
    assign rom[13'h0026] = 0;
    assign rom[13'h0027] = 0;
    assign rom[13'h0028] = 0;
    assign rom[13'h0029] = 0;
    assign rom[13'h002a] = 0;
    assign rom[13'h002b] = 0;
    assign rom[13'h002c] = 0;
    assign rom[13'h002d] = 0;
    assign rom[13'h002e] = 0;
    assign rom[13'h002f] = 0;
    assign rom[13'h0030] = 0;
    assign rom[13'h0031] = 0;
    assign rom[13'h0032] = 0;
    assign rom[13'h0033] = 0;
    assign rom[13'h0034] = 0;
    assign rom[13'h0035] = 0;
    assign rom[13'h0036] = 0;
    assign rom[13'h0037] = 0;
    assign rom[13'h0038] = 0;
    assign rom[13'h0039] = 0;
    assign rom[13'h003a] = 0;
    assign rom[13'h003b] = 0;
    assign rom[13'h003c] = 0;
    assign rom[13'h003d] = 0;
    assign rom[13'h003e] = 0;
    assign rom[13'h003f] = 0;
    assign rom[13'h0040] = 0;
    assign rom[13'h0041] = 0;
    assign rom[13'h0042] = 0;
    assign rom[13'h0043] = 0;
    assign rom[13'h0044] = 0;
    assign rom[13'h0045] = 0;
    assign rom[13'h0046] = 0;
    assign rom[13'h0047] = 0;
    assign rom[13'h0048] = 0;
    assign rom[13'h0049] = 0;
    assign rom[13'h004a] = 0;
    assign rom[13'h004b] = 0;
    assign rom[13'h004c] = 0;
    assign rom[13'h004d] = 0;
    assign rom[13'h004e] = 0;
    assign rom[13'h004f] = 0;
    assign rom[13'h0050] = 0;
    assign rom[13'h0051] = 0;
    assign rom[13'h0052] = 0;
    assign rom[13'h0053] = 0;
    assign rom[13'h0054] = 0;
    assign rom[13'h0055] = 0;
    assign rom[13'h0056] = 0;
    assign rom[13'h0057] = 0;
    assign rom[13'h0058] = 0;
    assign rom[13'h0059] = 0;
    assign rom[13'h005a] = 0;
    assign rom[13'h005b] = 0;
    assign rom[13'h005c] = 0;
    assign rom[13'h005d] = 0;
    assign rom[13'h005e] = 0;
    assign rom[13'h005f] = 0;
    assign rom[13'h0060] = 0;
    assign rom[13'h0061] = 0;
    assign rom[13'h0062] = 0;
    assign rom[13'h0063] = 0;
    assign rom[13'h0064] = 0;
    assign rom[13'h0065] = 0;
    assign rom[13'h0066] = 0;
    assign rom[13'h0067] = 0;
    assign rom[13'h0068] = 0;
    assign rom[13'h0069] = 0;
    assign rom[13'h006a] = 0;
    assign rom[13'h006b] = 0;
    assign rom[13'h006c] = 0;
    assign rom[13'h006d] = 0;
    assign rom[13'h006e] = 0;
    assign rom[13'h006f] = 0;
    assign rom[13'h0070] = 0;
    assign rom[13'h0071] = 0;
    assign rom[13'h0072] = 0;
    assign rom[13'h0073] = 0;
    assign rom[13'h0074] = 0;
    assign rom[13'h0075] = 0;
    assign rom[13'h0076] = 0;
    assign rom[13'h0077] = 0;
    assign rom[13'h0078] = 0;
    assign rom[13'h0079] = 0;
    assign rom[13'h007a] = 0;
    assign rom[13'h007b] = 0;
    assign rom[13'h007c] = 0;
    assign rom[13'h007d] = 0;
    assign rom[13'h007e] = 0;
    assign rom[13'h007f] = 0;
    assign rom[13'h0080] = 0;
    assign rom[13'h0081] = 0;
    assign rom[13'h0082] = 0;
    assign rom[13'h0083] = 0;
    assign rom[13'h0084] = 0;
    assign rom[13'h0085] = 0;
    assign rom[13'h0086] = 0;
    assign rom[13'h0087] = 0;
    assign rom[13'h0088] = 0;
    assign rom[13'h0089] = 0;
    assign rom[13'h008a] = 0;
    assign rom[13'h008b] = 0;
    assign rom[13'h008c] = 0;
    assign rom[13'h008d] = 0;
    assign rom[13'h008e] = 0;
    assign rom[13'h008f] = 0;
    assign rom[13'h0090] = 0;
    assign rom[13'h0091] = 0;
    assign rom[13'h0092] = 0;
    assign rom[13'h0093] = 0;
    assign rom[13'h0094] = 0;
    assign rom[13'h0095] = 0;
    assign rom[13'h0096] = 0;
    assign rom[13'h0097] = 0;
    assign rom[13'h0098] = 0;
    assign rom[13'h0099] = 0;
    assign rom[13'h009a] = 0;
    assign rom[13'h009b] = 0;
    assign rom[13'h009c] = 0;
    assign rom[13'h009d] = 0;
    assign rom[13'h009e] = 0;
    assign rom[13'h009f] = 0;
    assign rom[13'h00a0] = 0;
    assign rom[13'h00a1] = 0;
    assign rom[13'h00a2] = 0;
    assign rom[13'h00a3] = 0;
    assign rom[13'h00a4] = 0;
    assign rom[13'h00a5] = 0;
    assign rom[13'h00a6] = 0;
    assign rom[13'h00a7] = 0;
    assign rom[13'h00a8] = 0;
    assign rom[13'h00a9] = 0;
    assign rom[13'h00aa] = 0;
    assign rom[13'h00ab] = 0;
    assign rom[13'h00ac] = 0;
    assign rom[13'h00ad] = 0;
    assign rom[13'h00ae] = 0;
    assign rom[13'h00af] = 0;
    assign rom[13'h00b0] = 0;
    assign rom[13'h00b1] = 0;
    assign rom[13'h00b2] = 0;
    assign rom[13'h00b3] = 0;
    assign rom[13'h00b4] = 0;
    assign rom[13'h00b5] = 0;
    assign rom[13'h00b6] = 0;
    assign rom[13'h00b7] = 0;
    assign rom[13'h00b8] = 0;
    assign rom[13'h00b9] = 0;
    assign rom[13'h00ba] = 0;
    assign rom[13'h00bb] = 0;
    assign rom[13'h00bc] = 0;
    assign rom[13'h00bd] = 0;
    assign rom[13'h00be] = 0;
    assign rom[13'h00bf] = 0;
    assign rom[13'h00c0] = 0;
    assign rom[13'h00c1] = 0;
    assign rom[13'h00c2] = 0;
    assign rom[13'h00c3] = 0;
    assign rom[13'h00c4] = 0;
    assign rom[13'h00c5] = 0;
    assign rom[13'h00c6] = 0;
    assign rom[13'h00c7] = 0;
    assign rom[13'h00c8] = 0;
    assign rom[13'h00c9] = 0;
    assign rom[13'h00ca] = 0;
    assign rom[13'h00cb] = 0;
    assign rom[13'h00cc] = 0;
    assign rom[13'h00cd] = 0;
    assign rom[13'h00ce] = 0;
    assign rom[13'h00cf] = 0;
    assign rom[13'h00d0] = 0;
    assign rom[13'h00d1] = 0;
    assign rom[13'h00d2] = 0;
    assign rom[13'h00d3] = 0;
    assign rom[13'h00d4] = 0;
    assign rom[13'h00d5] = 0;
    assign rom[13'h00d6] = 0;
    assign rom[13'h00d7] = 0;
    assign rom[13'h00d8] = 0;
    assign rom[13'h00d9] = 0;
    assign rom[13'h00da] = 0;
    assign rom[13'h00db] = 0;
    assign rom[13'h00dc] = 0;
    assign rom[13'h00dd] = 0;
    assign rom[13'h00de] = 0;
    assign rom[13'h00df] = 0;
    assign rom[13'h00e0] = 0;
    assign rom[13'h00e1] = 0;
    assign rom[13'h00e2] = 0;
    assign rom[13'h00e3] = 0;
    assign rom[13'h00e4] = 0;
    assign rom[13'h00e5] = 0;
    assign rom[13'h00e6] = 0;
    assign rom[13'h00e7] = 0;
    assign rom[13'h00e8] = 0;
    assign rom[13'h00e9] = 0;
    assign rom[13'h00ea] = 0;
    assign rom[13'h00eb] = 0;
    assign rom[13'h00ec] = 0;
    assign rom[13'h00ed] = 0;
    assign rom[13'h00ee] = 0;
    assign rom[13'h00ef] = 0;
    assign rom[13'h00f0] = 0;
    assign rom[13'h00f1] = 0;
    assign rom[13'h00f2] = 0;
    assign rom[13'h00f3] = 0;
    assign rom[13'h00f4] = 0;
    assign rom[13'h00f5] = 0;
    assign rom[13'h00f6] = 0;
    assign rom[13'h00f7] = 0;
    assign rom[13'h00f8] = 0;
    assign rom[13'h00f9] = 0;
    assign rom[13'h00fa] = 0;
    assign rom[13'h00fb] = 0;
    assign rom[13'h00fc] = 0;
    assign rom[13'h00fd] = 0;
    assign rom[13'h00fe] = 0;
    assign rom[13'h00ff] = 0;
    assign rom[13'h0100] = 0;
    assign rom[13'h0101] = 0;
    assign rom[13'h0102] = 0;
    assign rom[13'h0103] = 0;
    assign rom[13'h0104] = 0;
    assign rom[13'h0105] = 0;
    assign rom[13'h0106] = 0;
    assign rom[13'h0107] = 0;
    assign rom[13'h0108] = 0;
    assign rom[13'h0109] = 0;
    assign rom[13'h010a] = 0;
    assign rom[13'h010b] = 0;
    assign rom[13'h010c] = 0;
    assign rom[13'h010d] = 0;
    assign rom[13'h010e] = 0;
    assign rom[13'h010f] = 0;
    assign rom[13'h0110] = 0;
    assign rom[13'h0111] = 0;
    assign rom[13'h0112] = 0;
    assign rom[13'h0113] = 0;
    assign rom[13'h0114] = 0;
    assign rom[13'h0115] = 0;
    assign rom[13'h0116] = 0;
    assign rom[13'h0117] = 0;
    assign rom[13'h0118] = 0;
    assign rom[13'h0119] = 0;
    assign rom[13'h011a] = 0;
    assign rom[13'h011b] = 0;
    assign rom[13'h011c] = 0;
    assign rom[13'h011d] = 0;
    assign rom[13'h011e] = 0;
    assign rom[13'h011f] = 0;
    assign rom[13'h0120] = 0;
    assign rom[13'h0121] = 0;
    assign rom[13'h0122] = 0;
    assign rom[13'h0123] = 0;
    assign rom[13'h0124] = 0;
    assign rom[13'h0125] = 0;
    assign rom[13'h0126] = 0;
    assign rom[13'h0127] = 0;
    assign rom[13'h0128] = 0;
    assign rom[13'h0129] = 0;
    assign rom[13'h012a] = 0;
    assign rom[13'h012b] = 0;
    assign rom[13'h012c] = 0;
    assign rom[13'h012d] = 0;
    assign rom[13'h012e] = 0;
    assign rom[13'h012f] = 0;
    assign rom[13'h0130] = 0;
    assign rom[13'h0131] = 0;
    assign rom[13'h0132] = 0;
    assign rom[13'h0133] = 0;
    assign rom[13'h0134] = 0;
    assign rom[13'h0135] = 0;
    assign rom[13'h0136] = 0;
    assign rom[13'h0137] = 0;
    assign rom[13'h0138] = 0;
    assign rom[13'h0139] = 0;
    assign rom[13'h013a] = 0;
    assign rom[13'h013b] = 0;
    assign rom[13'h013c] = 0;
    assign rom[13'h013d] = 0;
    assign rom[13'h013e] = 0;
    assign rom[13'h013f] = 0;
    assign rom[13'h0140] = 0;
    assign rom[13'h0141] = 0;
    assign rom[13'h0142] = 0;
    assign rom[13'h0143] = 0;
    assign rom[13'h0144] = 0;
    assign rom[13'h0145] = 0;
    assign rom[13'h0146] = 0;
    assign rom[13'h0147] = 0;
    assign rom[13'h0148] = 0;
    assign rom[13'h0149] = 0;
    assign rom[13'h014a] = 0;
    assign rom[13'h014b] = 0;
    assign rom[13'h014c] = 0;
    assign rom[13'h014d] = 0;
    assign rom[13'h014e] = 0;
    assign rom[13'h014f] = 0;
    assign rom[13'h0150] = 0;
    assign rom[13'h0151] = 0;
    assign rom[13'h0152] = 0;
    assign rom[13'h0153] = 0;
    assign rom[13'h0154] = 0;
    assign rom[13'h0155] = 0;
    assign rom[13'h0156] = 0;
    assign rom[13'h0157] = 0;
    assign rom[13'h0158] = 0;
    assign rom[13'h0159] = 0;
    assign rom[13'h015a] = 0;
    assign rom[13'h015b] = 0;
    assign rom[13'h015c] = 0;
    assign rom[13'h015d] = 0;
    assign rom[13'h015e] = 0;
    assign rom[13'h015f] = 0;
    assign rom[13'h0160] = 0;
    assign rom[13'h0161] = 0;
    assign rom[13'h0162] = 0;
    assign rom[13'h0163] = 0;
    assign rom[13'h0164] = 0;
    assign rom[13'h0165] = 0;
    assign rom[13'h0166] = 0;
    assign rom[13'h0167] = 0;
    assign rom[13'h0168] = 0;
    assign rom[13'h0169] = 0;
    assign rom[13'h016a] = 0;
    assign rom[13'h016b] = 0;
    assign rom[13'h016c] = 0;
    assign rom[13'h016d] = 0;
    assign rom[13'h016e] = 0;
    assign rom[13'h016f] = 0;
    assign rom[13'h0170] = 0;
    assign rom[13'h0171] = 0;
    assign rom[13'h0172] = 0;
    assign rom[13'h0173] = 0;
    assign rom[13'h0174] = 0;
    assign rom[13'h0175] = 0;
    assign rom[13'h0176] = 0;
    assign rom[13'h0177] = 0;
    assign rom[13'h0178] = 0;
    assign rom[13'h0179] = 0;
    assign rom[13'h017a] = 0;
    assign rom[13'h017b] = 0;
    assign rom[13'h017c] = 0;
    assign rom[13'h017d] = 0;
    assign rom[13'h017e] = 0;
    assign rom[13'h017f] = 0;
    assign rom[13'h0180] = 0;
    assign rom[13'h0181] = 0;
    assign rom[13'h0182] = 0;
    assign rom[13'h0183] = 0;
    assign rom[13'h0184] = 0;
    assign rom[13'h0185] = 0;
    assign rom[13'h0186] = 0;
    assign rom[13'h0187] = 0;
    assign rom[13'h0188] = 0;
    assign rom[13'h0189] = 0;
    assign rom[13'h018a] = 0;
    assign rom[13'h018b] = 0;
    assign rom[13'h018c] = 0;
    assign rom[13'h018d] = 0;
    assign rom[13'h018e] = 0;
    assign rom[13'h018f] = 0;
    assign rom[13'h0190] = 0;
    assign rom[13'h0191] = 0;
    assign rom[13'h0192] = 0;
    assign rom[13'h0193] = 0;
    assign rom[13'h0194] = 0;
    assign rom[13'h0195] = 0;
    assign rom[13'h0196] = 0;
    assign rom[13'h0197] = 0;
    assign rom[13'h0198] = 0;
    assign rom[13'h0199] = 0;
    assign rom[13'h019a] = 0;
    assign rom[13'h019b] = 0;
    assign rom[13'h019c] = 0;
    assign rom[13'h019d] = 0;
    assign rom[13'h019e] = 0;
    assign rom[13'h019f] = 0;
    assign rom[13'h01a0] = 0;
    assign rom[13'h01a1] = 0;
    assign rom[13'h01a2] = 0;
    assign rom[13'h01a3] = 0;
    assign rom[13'h01a4] = 0;
    assign rom[13'h01a5] = 0;
    assign rom[13'h01a6] = 0;
    assign rom[13'h01a7] = 0;
    assign rom[13'h01a8] = 0;
    assign rom[13'h01a9] = 0;
    assign rom[13'h01aa] = 0;
    assign rom[13'h01ab] = 0;
    assign rom[13'h01ac] = 0;
    assign rom[13'h01ad] = 0;
    assign rom[13'h01ae] = 0;
    assign rom[13'h01af] = 0;
    assign rom[13'h01b0] = 0;
    assign rom[13'h01b1] = 0;
    assign rom[13'h01b2] = 0;
    assign rom[13'h01b3] = 0;
    assign rom[13'h01b4] = 0;
    assign rom[13'h01b5] = 0;
    assign rom[13'h01b6] = 0;
    assign rom[13'h01b7] = 0;
    assign rom[13'h01b8] = 0;
    assign rom[13'h01b9] = 0;
    assign rom[13'h01ba] = 0;
    assign rom[13'h01bb] = 0;
    assign rom[13'h01bc] = 0;
    assign rom[13'h01bd] = 0;
    assign rom[13'h01be] = 0;
    assign rom[13'h01bf] = 0;
    assign rom[13'h01c0] = 0;
    assign rom[13'h01c1] = 0;
    assign rom[13'h01c2] = 0;
    assign rom[13'h01c3] = 0;
    assign rom[13'h01c4] = 0;
    assign rom[13'h01c5] = 0;
    assign rom[13'h01c6] = 0;
    assign rom[13'h01c7] = 0;
    assign rom[13'h01c8] = 0;
    assign rom[13'h01c9] = 0;
    assign rom[13'h01ca] = 0;
    assign rom[13'h01cb] = 0;
    assign rom[13'h01cc] = 0;
    assign rom[13'h01cd] = 0;
    assign rom[13'h01ce] = 0;
    assign rom[13'h01cf] = 0;
    assign rom[13'h01d0] = 0;
    assign rom[13'h01d1] = 0;
    assign rom[13'h01d2] = 0;
    assign rom[13'h01d3] = 0;
    assign rom[13'h01d4] = 0;
    assign rom[13'h01d5] = 0;
    assign rom[13'h01d6] = 0;
    assign rom[13'h01d7] = 0;
    assign rom[13'h01d8] = 0;
    assign rom[13'h01d9] = 0;
    assign rom[13'h01da] = 0;
    assign rom[13'h01db] = 0;
    assign rom[13'h01dc] = 0;
    assign rom[13'h01dd] = 0;
    assign rom[13'h01de] = 0;
    assign rom[13'h01df] = 0;
    assign rom[13'h01e0] = 0;
    assign rom[13'h01e1] = 0;
    assign rom[13'h01e2] = 0;
    assign rom[13'h01e3] = 0;
    assign rom[13'h01e4] = 0;
    assign rom[13'h01e5] = 0;
    assign rom[13'h01e6] = 0;
    assign rom[13'h01e7] = 0;
    assign rom[13'h01e8] = 0;
    assign rom[13'h01e9] = 0;
    assign rom[13'h01ea] = 0;
    assign rom[13'h01eb] = 0;
    assign rom[13'h01ec] = 0;
    assign rom[13'h01ed] = 0;
    assign rom[13'h01ee] = 0;
    assign rom[13'h01ef] = 0;
    assign rom[13'h01f0] = 0;
    assign rom[13'h01f1] = 0;
    assign rom[13'h01f2] = 0;
    assign rom[13'h01f3] = 0;
    assign rom[13'h01f4] = 0;
    assign rom[13'h01f5] = 0;
    assign rom[13'h01f6] = 0;
    assign rom[13'h01f7] = 0;
    assign rom[13'h01f8] = 0;
    assign rom[13'h01f9] = 0;
    assign rom[13'h01fa] = 0;
    assign rom[13'h01fb] = 0;
    assign rom[13'h01fc] = 0;
    assign rom[13'h01fd] = 0;
    assign rom[13'h01fe] = 0;
    assign rom[13'h01ff] = 0;
    assign rom[13'h0200] = 0;
    assign rom[13'h0201] = 0;
    assign rom[13'h0202] = 0;
    assign rom[13'h0203] = 0;
    assign rom[13'h0204] = 0;
    assign rom[13'h0205] = 0;
    assign rom[13'h0206] = 0;
    assign rom[13'h0207] = 0;
    assign rom[13'h0208] = 0;
    assign rom[13'h0209] = 0;
    assign rom[13'h020a] = 0;
    assign rom[13'h020b] = 0;
    assign rom[13'h020c] = 0;
    assign rom[13'h020d] = 0;
    assign rom[13'h020e] = 0;
    assign rom[13'h020f] = 0;
    assign rom[13'h0210] = 0;
    assign rom[13'h0211] = 0;
    assign rom[13'h0212] = 0;
    assign rom[13'h0213] = 0;
    assign rom[13'h0214] = 0;
    assign rom[13'h0215] = 0;
    assign rom[13'h0216] = 0;
    assign rom[13'h0217] = 0;
    assign rom[13'h0218] = 0;
    assign rom[13'h0219] = 0;
    assign rom[13'h021a] = 0;
    assign rom[13'h021b] = 0;
    assign rom[13'h021c] = 0;
    assign rom[13'h021d] = 0;
    assign rom[13'h021e] = 0;
    assign rom[13'h021f] = 0;
    assign rom[13'h0220] = 0;
    assign rom[13'h0221] = 0;
    assign rom[13'h0222] = 0;
    assign rom[13'h0223] = 0;
    assign rom[13'h0224] = 0;
    assign rom[13'h0225] = 0;
    assign rom[13'h0226] = 0;
    assign rom[13'h0227] = 0;
    assign rom[13'h0228] = 0;
    assign rom[13'h0229] = 0;
    assign rom[13'h022a] = 0;
    assign rom[13'h022b] = 0;
    assign rom[13'h022c] = 0;
    assign rom[13'h022d] = 0;
    assign rom[13'h022e] = 0;
    assign rom[13'h022f] = 0;
    assign rom[13'h0230] = 0;
    assign rom[13'h0231] = 0;
    assign rom[13'h0232] = 0;
    assign rom[13'h0233] = 0;
    assign rom[13'h0234] = 0;
    assign rom[13'h0235] = 0;
    assign rom[13'h0236] = 0;
    assign rom[13'h0237] = 0;
    assign rom[13'h0238] = 0;
    assign rom[13'h0239] = 0;
    assign rom[13'h023a] = 0;
    assign rom[13'h023b] = 0;
    assign rom[13'h023c] = 0;
    assign rom[13'h023d] = 0;
    assign rom[13'h023e] = 0;
    assign rom[13'h023f] = 0;
    assign rom[13'h0240] = 0;
    assign rom[13'h0241] = 0;
    assign rom[13'h0242] = 0;
    assign rom[13'h0243] = 0;
    assign rom[13'h0244] = 0;
    assign rom[13'h0245] = 0;
    assign rom[13'h0246] = 0;
    assign rom[13'h0247] = 0;
    assign rom[13'h0248] = 0;
    assign rom[13'h0249] = 0;
    assign rom[13'h024a] = 0;
    assign rom[13'h024b] = 0;
    assign rom[13'h024c] = 0;
    assign rom[13'h024d] = 0;
    assign rom[13'h024e] = 0;
    assign rom[13'h024f] = 0;
    assign rom[13'h0250] = 0;
    assign rom[13'h0251] = 0;
    assign rom[13'h0252] = 0;
    assign rom[13'h0253] = 0;
    assign rom[13'h0254] = 0;
    assign rom[13'h0255] = 0;
    assign rom[13'h0256] = 0;
    assign rom[13'h0257] = 0;
    assign rom[13'h0258] = 0;
    assign rom[13'h0259] = 0;
    assign rom[13'h025a] = 0;
    assign rom[13'h025b] = 0;
    assign rom[13'h025c] = 0;
    assign rom[13'h025d] = 0;
    assign rom[13'h025e] = 0;
    assign rom[13'h025f] = 0;
    assign rom[13'h0260] = 0;
    assign rom[13'h0261] = 0;
    assign rom[13'h0262] = 0;
    assign rom[13'h0263] = 0;
    assign rom[13'h0264] = 0;
    assign rom[13'h0265] = 0;
    assign rom[13'h0266] = 0;
    assign rom[13'h0267] = 0;
    assign rom[13'h0268] = 0;
    assign rom[13'h0269] = 0;
    assign rom[13'h026a] = 0;
    assign rom[13'h026b] = 0;
    assign rom[13'h026c] = 0;
    assign rom[13'h026d] = 0;
    assign rom[13'h026e] = 0;
    assign rom[13'h026f] = 0;
    assign rom[13'h0270] = 0;
    assign rom[13'h0271] = 0;
    assign rom[13'h0272] = 0;
    assign rom[13'h0273] = 0;
    assign rom[13'h0274] = 0;
    assign rom[13'h0275] = 0;
    assign rom[13'h0276] = 0;
    assign rom[13'h0277] = 0;
    assign rom[13'h0278] = 0;
    assign rom[13'h0279] = 0;
    assign rom[13'h027a] = 0;
    assign rom[13'h027b] = 0;
    assign rom[13'h027c] = 0;
    assign rom[13'h027d] = 0;
    assign rom[13'h027e] = 0;
    assign rom[13'h027f] = 0;
    assign rom[13'h0280] = 0;
    assign rom[13'h0281] = 0;
    assign rom[13'h0282] = 0;
    assign rom[13'h0283] = 0;
    assign rom[13'h0284] = 0;
    assign rom[13'h0285] = 0;
    assign rom[13'h0286] = 0;
    assign rom[13'h0287] = 0;
    assign rom[13'h0288] = 0;
    assign rom[13'h0289] = 0;
    assign rom[13'h028a] = 0;
    assign rom[13'h028b] = 0;
    assign rom[13'h028c] = 0;
    assign rom[13'h028d] = 0;
    assign rom[13'h028e] = 0;
    assign rom[13'h028f] = 0;
    assign rom[13'h0290] = 0;
    assign rom[13'h0291] = 0;
    assign rom[13'h0292] = 0;
    assign rom[13'h0293] = 0;
    assign rom[13'h0294] = 0;
    assign rom[13'h0295] = 0;
    assign rom[13'h0296] = 0;
    assign rom[13'h0297] = 0;
    assign rom[13'h0298] = 0;
    assign rom[13'h0299] = 0;
    assign rom[13'h029a] = 0;
    assign rom[13'h029b] = 0;
    assign rom[13'h029c] = 0;
    assign rom[13'h029d] = 0;
    assign rom[13'h029e] = 0;
    assign rom[13'h029f] = 0;
    assign rom[13'h02a0] = 0;
    assign rom[13'h02a1] = 0;
    assign rom[13'h02a2] = 0;
    assign rom[13'h02a3] = 0;
    assign rom[13'h02a4] = 0;
    assign rom[13'h02a5] = 0;
    assign rom[13'h02a6] = 0;
    assign rom[13'h02a7] = 0;
    assign rom[13'h02a8] = 0;
    assign rom[13'h02a9] = 0;
    assign rom[13'h02aa] = 0;
    assign rom[13'h02ab] = 0;
    assign rom[13'h02ac] = 0;
    assign rom[13'h02ad] = 0;
    assign rom[13'h02ae] = 0;
    assign rom[13'h02af] = 0;
    assign rom[13'h02b0] = 0;
    assign rom[13'h02b1] = 0;
    assign rom[13'h02b2] = 0;
    assign rom[13'h02b3] = 0;
    assign rom[13'h02b4] = 0;
    assign rom[13'h02b5] = 0;
    assign rom[13'h02b6] = 0;
    assign rom[13'h02b7] = 0;
    assign rom[13'h02b8] = 0;
    assign rom[13'h02b9] = 0;
    assign rom[13'h02ba] = 0;
    assign rom[13'h02bb] = 0;
    assign rom[13'h02bc] = 0;
    assign rom[13'h02bd] = 0;
    assign rom[13'h02be] = 0;
    assign rom[13'h02bf] = 0;
    assign rom[13'h02c0] = 0;
    assign rom[13'h02c1] = 0;
    assign rom[13'h02c2] = 0;
    assign rom[13'h02c3] = 0;
    assign rom[13'h02c4] = 0;
    assign rom[13'h02c5] = 0;
    assign rom[13'h02c6] = 0;
    assign rom[13'h02c7] = 0;
    assign rom[13'h02c8] = 0;
    assign rom[13'h02c9] = 0;
    assign rom[13'h02ca] = 0;
    assign rom[13'h02cb] = 0;
    assign rom[13'h02cc] = 0;
    assign rom[13'h02cd] = 0;
    assign rom[13'h02ce] = 0;
    assign rom[13'h02cf] = 0;
    assign rom[13'h02d0] = 0;
    assign rom[13'h02d1] = 0;
    assign rom[13'h02d2] = 0;
    assign rom[13'h02d3] = 0;
    assign rom[13'h02d4] = 0;
    assign rom[13'h02d5] = 0;
    assign rom[13'h02d6] = 0;
    assign rom[13'h02d7] = 0;
    assign rom[13'h02d8] = 0;
    assign rom[13'h02d9] = 0;
    assign rom[13'h02da] = 0;
    assign rom[13'h02db] = 0;
    assign rom[13'h02dc] = 0;
    assign rom[13'h02dd] = 0;
    assign rom[13'h02de] = 0;
    assign rom[13'h02df] = 0;
    assign rom[13'h02e0] = 0;
    assign rom[13'h02e1] = 0;
    assign rom[13'h02e2] = 0;
    assign rom[13'h02e3] = 0;
    assign rom[13'h02e4] = 0;
    assign rom[13'h02e5] = 0;
    assign rom[13'h02e6] = 0;
    assign rom[13'h02e7] = 0;
    assign rom[13'h02e8] = 0;
    assign rom[13'h02e9] = 0;
    assign rom[13'h02ea] = 0;
    assign rom[13'h02eb] = 0;
    assign rom[13'h02ec] = 0;
    assign rom[13'h02ed] = 0;
    assign rom[13'h02ee] = 0;
    assign rom[13'h02ef] = 0;
    assign rom[13'h02f0] = 0;
    assign rom[13'h02f1] = 0;
    assign rom[13'h02f2] = 0;
    assign rom[13'h02f3] = 0;
    assign rom[13'h02f4] = 0;
    assign rom[13'h02f5] = 0;
    assign rom[13'h02f6] = 0;
    assign rom[13'h02f7] = 0;
    assign rom[13'h02f8] = 0;
    assign rom[13'h02f9] = 0;
    assign rom[13'h02fa] = 0;
    assign rom[13'h02fb] = 0;
    assign rom[13'h02fc] = 0;
    assign rom[13'h02fd] = 0;
    assign rom[13'h02fe] = 0;
    assign rom[13'h02ff] = 0;
    assign rom[13'h0300] = 0;
    assign rom[13'h0301] = 0;
    assign rom[13'h0302] = 0;
    assign rom[13'h0303] = 0;
    assign rom[13'h0304] = 0;
    assign rom[13'h0305] = 0;
    assign rom[13'h0306] = 0;
    assign rom[13'h0307] = 0;
    assign rom[13'h0308] = 0;
    assign rom[13'h0309] = 0;
    assign rom[13'h030a] = 0;
    assign rom[13'h030b] = 0;
    assign rom[13'h030c] = 0;
    assign rom[13'h030d] = 0;
    assign rom[13'h030e] = 0;
    assign rom[13'h030f] = 0;
    assign rom[13'h0310] = 0;
    assign rom[13'h0311] = 0;
    assign rom[13'h0312] = 0;
    assign rom[13'h0313] = 0;
    assign rom[13'h0314] = 0;
    assign rom[13'h0315] = 0;
    assign rom[13'h0316] = 0;
    assign rom[13'h0317] = 0;
    assign rom[13'h0318] = 0;
    assign rom[13'h0319] = 0;
    assign rom[13'h031a] = 0;
    assign rom[13'h031b] = 0;
    assign rom[13'h031c] = 0;
    assign rom[13'h031d] = 0;
    assign rom[13'h031e] = 0;
    assign rom[13'h031f] = 0;
    assign rom[13'h0320] = 0;
    assign rom[13'h0321] = 0;
    assign rom[13'h0322] = 0;
    assign rom[13'h0323] = 0;
    assign rom[13'h0324] = 0;
    assign rom[13'h0325] = 0;
    assign rom[13'h0326] = 0;
    assign rom[13'h0327] = 0;
    assign rom[13'h0328] = 0;
    assign rom[13'h0329] = 0;
    assign rom[13'h032a] = 0;
    assign rom[13'h032b] = 0;
    assign rom[13'h032c] = 0;
    assign rom[13'h032d] = 0;
    assign rom[13'h032e] = 0;
    assign rom[13'h032f] = 0;
    assign rom[13'h0330] = 0;
    assign rom[13'h0331] = 0;
    assign rom[13'h0332] = 0;
    assign rom[13'h0333] = 0;
    assign rom[13'h0334] = 0;
    assign rom[13'h0335] = 0;
    assign rom[13'h0336] = 0;
    assign rom[13'h0337] = 0;
    assign rom[13'h0338] = 0;
    assign rom[13'h0339] = 0;
    assign rom[13'h033a] = 0;
    assign rom[13'h033b] = 0;
    assign rom[13'h033c] = 0;
    assign rom[13'h033d] = 0;
    assign rom[13'h033e] = 0;
    assign rom[13'h033f] = 0;
    assign rom[13'h0340] = 0;
    assign rom[13'h0341] = 0;
    assign rom[13'h0342] = 0;
    assign rom[13'h0343] = 0;
    assign rom[13'h0344] = 0;
    assign rom[13'h0345] = 0;
    assign rom[13'h0346] = 0;
    assign rom[13'h0347] = 0;
    assign rom[13'h0348] = 0;
    assign rom[13'h0349] = 0;
    assign rom[13'h034a] = 0;
    assign rom[13'h034b] = 0;
    assign rom[13'h034c] = 0;
    assign rom[13'h034d] = 0;
    assign rom[13'h034e] = 0;
    assign rom[13'h034f] = 0;
    assign rom[13'h0350] = 0;
    assign rom[13'h0351] = 0;
    assign rom[13'h0352] = 0;
    assign rom[13'h0353] = 0;
    assign rom[13'h0354] = 0;
    assign rom[13'h0355] = 0;
    assign rom[13'h0356] = 0;
    assign rom[13'h0357] = 0;
    assign rom[13'h0358] = 0;
    assign rom[13'h0359] = 0;
    assign rom[13'h035a] = 0;
    assign rom[13'h035b] = 0;
    assign rom[13'h035c] = 0;
    assign rom[13'h035d] = 0;
    assign rom[13'h035e] = 0;
    assign rom[13'h035f] = 0;
    assign rom[13'h0360] = 0;
    assign rom[13'h0361] = 0;
    assign rom[13'h0362] = 0;
    assign rom[13'h0363] = 0;
    assign rom[13'h0364] = 0;
    assign rom[13'h0365] = 0;
    assign rom[13'h0366] = 0;
    assign rom[13'h0367] = 0;
    assign rom[13'h0368] = 0;
    assign rom[13'h0369] = 0;
    assign rom[13'h036a] = 0;
    assign rom[13'h036b] = 0;
    assign rom[13'h036c] = 0;
    assign rom[13'h036d] = 0;
    assign rom[13'h036e] = 0;
    assign rom[13'h036f] = 0;
    assign rom[13'h0370] = 0;
    assign rom[13'h0371] = 0;
    assign rom[13'h0372] = 0;
    assign rom[13'h0373] = 0;
    assign rom[13'h0374] = 0;
    assign rom[13'h0375] = 0;
    assign rom[13'h0376] = 0;
    assign rom[13'h0377] = 0;
    assign rom[13'h0378] = 0;
    assign rom[13'h0379] = 0;
    assign rom[13'h037a] = 0;
    assign rom[13'h037b] = 0;
    assign rom[13'h037c] = 0;
    assign rom[13'h037d] = 0;
    assign rom[13'h037e] = 0;
    assign rom[13'h037f] = 0;
    assign rom[13'h0380] = 0;
    assign rom[13'h0381] = 0;
    assign rom[13'h0382] = 0;
    assign rom[13'h0383] = 0;
    assign rom[13'h0384] = 0;
    assign rom[13'h0385] = 0;
    assign rom[13'h0386] = 0;
    assign rom[13'h0387] = 0;
    assign rom[13'h0388] = 0;
    assign rom[13'h0389] = 0;
    assign rom[13'h038a] = 0;
    assign rom[13'h038b] = 0;
    assign rom[13'h038c] = 0;
    assign rom[13'h038d] = 0;
    assign rom[13'h038e] = 0;
    assign rom[13'h038f] = 0;
    assign rom[13'h0390] = 0;
    assign rom[13'h0391] = 0;
    assign rom[13'h0392] = 0;
    assign rom[13'h0393] = 0;
    assign rom[13'h0394] = 0;
    assign rom[13'h0395] = 0;
    assign rom[13'h0396] = 0;
    assign rom[13'h0397] = 0;
    assign rom[13'h0398] = 0;
    assign rom[13'h0399] = 0;
    assign rom[13'h039a] = 0;
    assign rom[13'h039b] = 0;
    assign rom[13'h039c] = 0;
    assign rom[13'h039d] = 0;
    assign rom[13'h039e] = 0;
    assign rom[13'h039f] = 0;
    assign rom[13'h03a0] = 0;
    assign rom[13'h03a1] = 0;
    assign rom[13'h03a2] = 0;
    assign rom[13'h03a3] = 0;
    assign rom[13'h03a4] = 0;
    assign rom[13'h03a5] = 0;
    assign rom[13'h03a6] = 0;
    assign rom[13'h03a7] = 0;
    assign rom[13'h03a8] = 0;
    assign rom[13'h03a9] = 0;
    assign rom[13'h03aa] = 0;
    assign rom[13'h03ab] = 0;
    assign rom[13'h03ac] = 0;
    assign rom[13'h03ad] = 0;
    assign rom[13'h03ae] = 0;
    assign rom[13'h03af] = 0;
    assign rom[13'h03b0] = 0;
    assign rom[13'h03b1] = 0;
    assign rom[13'h03b2] = 0;
    assign rom[13'h03b3] = 0;
    assign rom[13'h03b4] = 0;
    assign rom[13'h03b5] = 0;
    assign rom[13'h03b6] = 0;
    assign rom[13'h03b7] = 0;
    assign rom[13'h03b8] = 0;
    assign rom[13'h03b9] = 0;
    assign rom[13'h03ba] = 0;
    assign rom[13'h03bb] = 0;
    assign rom[13'h03bc] = 0;
    assign rom[13'h03bd] = 0;
    assign rom[13'h03be] = 0;
    assign rom[13'h03bf] = 0;
    assign rom[13'h03c0] = 0;
    assign rom[13'h03c1] = 0;
    assign rom[13'h03c2] = 0;
    assign rom[13'h03c3] = 0;
    assign rom[13'h03c4] = 0;
    assign rom[13'h03c5] = 0;
    assign rom[13'h03c6] = 0;
    assign rom[13'h03c7] = 0;
    assign rom[13'h03c8] = 0;
    assign rom[13'h03c9] = 0;
    assign rom[13'h03ca] = 0;
    assign rom[13'h03cb] = 0;
    assign rom[13'h03cc] = 0;
    assign rom[13'h03cd] = 0;
    assign rom[13'h03ce] = 0;
    assign rom[13'h03cf] = 0;
    assign rom[13'h03d0] = 0;
    assign rom[13'h03d1] = 0;
    assign rom[13'h03d2] = 0;
    assign rom[13'h03d3] = 0;
    assign rom[13'h03d4] = 0;
    assign rom[13'h03d5] = 0;
    assign rom[13'h03d6] = 0;
    assign rom[13'h03d7] = 0;
    assign rom[13'h03d8] = 0;
    assign rom[13'h03d9] = 0;
    assign rom[13'h03da] = 0;
    assign rom[13'h03db] = 0;
    assign rom[13'h03dc] = 0;
    assign rom[13'h03dd] = 0;
    assign rom[13'h03de] = 0;
    assign rom[13'h03df] = 0;
    assign rom[13'h03e0] = 0;
    assign rom[13'h03e1] = 0;
    assign rom[13'h03e2] = 0;
    assign rom[13'h03e3] = 0;
    assign rom[13'h03e4] = 0;
    assign rom[13'h03e5] = 0;
    assign rom[13'h03e6] = 0;
    assign rom[13'h03e7] = 0;
    assign rom[13'h03e8] = 0;
    assign rom[13'h03e9] = 0;
    assign rom[13'h03ea] = 0;
    assign rom[13'h03eb] = 0;
    assign rom[13'h03ec] = 0;
    assign rom[13'h03ed] = 0;
    assign rom[13'h03ee] = 0;
    assign rom[13'h03ef] = 0;
    assign rom[13'h03f0] = 0;
    assign rom[13'h03f1] = 0;
    assign rom[13'h03f2] = 0;
    assign rom[13'h03f3] = 0;
    assign rom[13'h03f4] = 0;
    assign rom[13'h03f5] = 0;
    assign rom[13'h03f6] = 0;
    assign rom[13'h03f7] = 0;
    assign rom[13'h03f8] = 0;
    assign rom[13'h03f9] = 0;
    assign rom[13'h03fa] = 0;
    assign rom[13'h03fb] = 0;
    assign rom[13'h03fc] = 0;
    assign rom[13'h03fd] = 0;
    assign rom[13'h03fe] = 0;
    assign rom[13'h03ff] = 0;
    assign rom[13'h0400] = 0;
    assign rom[13'h0401] = 0;
    assign rom[13'h0402] = 0;
    assign rom[13'h0403] = 0;
    assign rom[13'h0404] = 0;
    assign rom[13'h0405] = 0;
    assign rom[13'h0406] = 0;
    assign rom[13'h0407] = 0;
    assign rom[13'h0408] = 0;
    assign rom[13'h0409] = 0;
    assign rom[13'h040a] = 0;
    assign rom[13'h040b] = 0;
    assign rom[13'h040c] = 0;
    assign rom[13'h040d] = 0;
    assign rom[13'h040e] = 0;
    assign rom[13'h040f] = 0;
    assign rom[13'h0410] = 0;
    assign rom[13'h0411] = 0;
    assign rom[13'h0412] = 0;
    assign rom[13'h0413] = 0;
    assign rom[13'h0414] = 0;
    assign rom[13'h0415] = 0;
    assign rom[13'h0416] = 0;
    assign rom[13'h0417] = 0;
    assign rom[13'h0418] = 0;
    assign rom[13'h0419] = 0;
    assign rom[13'h041a] = 0;
    assign rom[13'h041b] = 0;
    assign rom[13'h041c] = 0;
    assign rom[13'h041d] = 0;
    assign rom[13'h041e] = 0;
    assign rom[13'h041f] = 0;
    assign rom[13'h0420] = 0;
    assign rom[13'h0421] = 0;
    assign rom[13'h0422] = 0;
    assign rom[13'h0423] = 0;
    assign rom[13'h0424] = 0;
    assign rom[13'h0425] = 0;
    assign rom[13'h0426] = 0;
    assign rom[13'h0427] = 0;
    assign rom[13'h0428] = 0;
    assign rom[13'h0429] = 0;
    assign rom[13'h042a] = 0;
    assign rom[13'h042b] = 0;
    assign rom[13'h042c] = 0;
    assign rom[13'h042d] = 0;
    assign rom[13'h042e] = 0;
    assign rom[13'h042f] = 0;
    assign rom[13'h0430] = 0;
    assign rom[13'h0431] = 0;
    assign rom[13'h0432] = 0;
    assign rom[13'h0433] = 0;
    assign rom[13'h0434] = 0;
    assign rom[13'h0435] = 0;
    assign rom[13'h0436] = 0;
    assign rom[13'h0437] = 0;
    assign rom[13'h0438] = 0;
    assign rom[13'h0439] = 0;
    assign rom[13'h043a] = 0;
    assign rom[13'h043b] = 0;
    assign rom[13'h043c] = 0;
    assign rom[13'h043d] = 0;
    assign rom[13'h043e] = 0;
    assign rom[13'h043f] = 0;
    assign rom[13'h0440] = 0;
    assign rom[13'h0441] = 0;
    assign rom[13'h0442] = 0;
    assign rom[13'h0443] = 0;
    assign rom[13'h0444] = 0;
    assign rom[13'h0445] = 0;
    assign rom[13'h0446] = 0;
    assign rom[13'h0447] = 0;
    assign rom[13'h0448] = 0;
    assign rom[13'h0449] = 0;
    assign rom[13'h044a] = 0;
    assign rom[13'h044b] = 0;
    assign rom[13'h044c] = 0;
    assign rom[13'h044d] = 0;
    assign rom[13'h044e] = 0;
    assign rom[13'h044f] = 0;
    assign rom[13'h0450] = 0;
    assign rom[13'h0451] = 0;
    assign rom[13'h0452] = 0;
    assign rom[13'h0453] = 0;
    assign rom[13'h0454] = 0;
    assign rom[13'h0455] = 0;
    assign rom[13'h0456] = 0;
    assign rom[13'h0457] = 0;
    assign rom[13'h0458] = 0;
    assign rom[13'h0459] = 0;
    assign rom[13'h045a] = 0;
    assign rom[13'h045b] = 0;
    assign rom[13'h045c] = 0;
    assign rom[13'h045d] = 0;
    assign rom[13'h045e] = 0;
    assign rom[13'h045f] = 0;
    assign rom[13'h0460] = 0;
    assign rom[13'h0461] = 0;
    assign rom[13'h0462] = 0;
    assign rom[13'h0463] = 0;
    assign rom[13'h0464] = 0;
    assign rom[13'h0465] = 0;
    assign rom[13'h0466] = 0;
    assign rom[13'h0467] = 0;
    assign rom[13'h0468] = 0;
    assign rom[13'h0469] = 0;
    assign rom[13'h046a] = 0;
    assign rom[13'h046b] = 0;
    assign rom[13'h046c] = 0;
    assign rom[13'h046d] = 0;
    assign rom[13'h046e] = 0;
    assign rom[13'h046f] = 0;
    assign rom[13'h0470] = 0;
    assign rom[13'h0471] = 0;
    assign rom[13'h0472] = 0;
    assign rom[13'h0473] = 0;
    assign rom[13'h0474] = 0;
    assign rom[13'h0475] = 0;
    assign rom[13'h0476] = 0;
    assign rom[13'h0477] = 0;
    assign rom[13'h0478] = 0;
    assign rom[13'h0479] = 0;
    assign rom[13'h047a] = 0;
    assign rom[13'h047b] = 0;
    assign rom[13'h047c] = 0;
    assign rom[13'h047d] = 0;
    assign rom[13'h047e] = 0;
    assign rom[13'h047f] = 0;
    assign rom[13'h0480] = 0;
    assign rom[13'h0481] = 0;
    assign rom[13'h0482] = 0;
    assign rom[13'h0483] = 0;
    assign rom[13'h0484] = 0;
    assign rom[13'h0485] = 0;
    assign rom[13'h0486] = 0;
    assign rom[13'h0487] = 0;
    assign rom[13'h0488] = 0;
    assign rom[13'h0489] = 0;
    assign rom[13'h048a] = 0;
    assign rom[13'h048b] = 0;
    assign rom[13'h048c] = 0;
    assign rom[13'h048d] = 0;
    assign rom[13'h048e] = 0;
    assign rom[13'h048f] = 0;
    assign rom[13'h0490] = 0;
    assign rom[13'h0491] = 0;
    assign rom[13'h0492] = 0;
    assign rom[13'h0493] = 0;
    assign rom[13'h0494] = 0;
    assign rom[13'h0495] = 0;
    assign rom[13'h0496] = 0;
    assign rom[13'h0497] = 0;
    assign rom[13'h0498] = 0;
    assign rom[13'h0499] = 0;
    assign rom[13'h049a] = 0;
    assign rom[13'h049b] = 0;
    assign rom[13'h049c] = 0;
    assign rom[13'h049d] = 0;
    assign rom[13'h049e] = 0;
    assign rom[13'h049f] = 0;
    assign rom[13'h04a0] = 0;
    assign rom[13'h04a1] = 0;
    assign rom[13'h04a2] = 0;
    assign rom[13'h04a3] = 0;
    assign rom[13'h04a4] = 0;
    assign rom[13'h04a5] = 0;
    assign rom[13'h04a6] = 0;
    assign rom[13'h04a7] = 0;
    assign rom[13'h04a8] = 0;
    assign rom[13'h04a9] = 0;
    assign rom[13'h04aa] = 0;
    assign rom[13'h04ab] = 0;
    assign rom[13'h04ac] = 0;
    assign rom[13'h04ad] = 0;
    assign rom[13'h04ae] = 0;
    assign rom[13'h04af] = 0;
    assign rom[13'h04b0] = 0;
    assign rom[13'h04b1] = 0;
    assign rom[13'h04b2] = 0;
    assign rom[13'h04b3] = 0;
    assign rom[13'h04b4] = 0;
    assign rom[13'h04b5] = 0;
    assign rom[13'h04b6] = 0;
    assign rom[13'h04b7] = 0;
    assign rom[13'h04b8] = 0;
    assign rom[13'h04b9] = 0;
    assign rom[13'h04ba] = 0;
    assign rom[13'h04bb] = 0;
    assign rom[13'h04bc] = 0;
    assign rom[13'h04bd] = 0;
    assign rom[13'h04be] = 0;
    assign rom[13'h04bf] = 0;
    assign rom[13'h04c0] = 0;
    assign rom[13'h04c1] = 0;
    assign rom[13'h04c2] = 0;
    assign rom[13'h04c3] = 0;
    assign rom[13'h04c4] = 0;
    assign rom[13'h04c5] = 0;
    assign rom[13'h04c6] = 0;
    assign rom[13'h04c7] = 0;
    assign rom[13'h04c8] = 0;
    assign rom[13'h04c9] = 0;
    assign rom[13'h04ca] = 0;
    assign rom[13'h04cb] = 0;
    assign rom[13'h04cc] = 0;
    assign rom[13'h04cd] = 0;
    assign rom[13'h04ce] = 0;
    assign rom[13'h04cf] = 0;
    assign rom[13'h04d0] = 0;
    assign rom[13'h04d1] = 0;
    assign rom[13'h04d2] = 0;
    assign rom[13'h04d3] = 0;
    assign rom[13'h04d4] = 0;
    assign rom[13'h04d5] = 0;
    assign rom[13'h04d6] = 0;
    assign rom[13'h04d7] = 0;
    assign rom[13'h04d8] = 0;
    assign rom[13'h04d9] = 0;
    assign rom[13'h04da] = 0;
    assign rom[13'h04db] = 0;
    assign rom[13'h04dc] = 0;
    assign rom[13'h04dd] = 0;
    assign rom[13'h04de] = 0;
    assign rom[13'h04df] = 0;
    assign rom[13'h04e0] = 0;
    assign rom[13'h04e1] = 0;
    assign rom[13'h04e2] = 0;
    assign rom[13'h04e3] = 0;
    assign rom[13'h04e4] = 0;
    assign rom[13'h04e5] = 0;
    assign rom[13'h04e6] = 0;
    assign rom[13'h04e7] = 0;
    assign rom[13'h04e8] = 0;
    assign rom[13'h04e9] = 0;
    assign rom[13'h04ea] = 0;
    assign rom[13'h04eb] = 0;
    assign rom[13'h04ec] = 0;
    assign rom[13'h04ed] = 0;
    assign rom[13'h04ee] = 0;
    assign rom[13'h04ef] = 0;
    assign rom[13'h04f0] = 0;
    assign rom[13'h04f1] = 0;
    assign rom[13'h04f2] = 0;
    assign rom[13'h04f3] = 0;
    assign rom[13'h04f4] = 0;
    assign rom[13'h04f5] = 0;
    assign rom[13'h04f6] = 0;
    assign rom[13'h04f7] = 0;
    assign rom[13'h04f8] = 0;
    assign rom[13'h04f9] = 0;
    assign rom[13'h04fa] = 0;
    assign rom[13'h04fb] = 0;
    assign rom[13'h04fc] = 0;
    assign rom[13'h04fd] = 0;
    assign rom[13'h04fe] = 0;
    assign rom[13'h04ff] = 0;
    assign rom[13'h0500] = 0;
    assign rom[13'h0501] = 0;
    assign rom[13'h0502] = 0;
    assign rom[13'h0503] = 0;
    assign rom[13'h0504] = 0;
    assign rom[13'h0505] = 0;
    assign rom[13'h0506] = 0;
    assign rom[13'h0507] = 0;
    assign rom[13'h0508] = 0;
    assign rom[13'h0509] = 0;
    assign rom[13'h050a] = 0;
    assign rom[13'h050b] = 0;
    assign rom[13'h050c] = 0;
    assign rom[13'h050d] = 0;
    assign rom[13'h050e] = 0;
    assign rom[13'h050f] = 0;
    assign rom[13'h0510] = 0;
    assign rom[13'h0511] = 0;
    assign rom[13'h0512] = 0;
    assign rom[13'h0513] = 0;
    assign rom[13'h0514] = 0;
    assign rom[13'h0515] = 0;
    assign rom[13'h0516] = 0;
    assign rom[13'h0517] = 0;
    assign rom[13'h0518] = 0;
    assign rom[13'h0519] = 0;
    assign rom[13'h051a] = 0;
    assign rom[13'h051b] = 0;
    assign rom[13'h051c] = 0;
    assign rom[13'h051d] = 0;
    assign rom[13'h051e] = 0;
    assign rom[13'h051f] = 0;
    assign rom[13'h0520] = 0;
    assign rom[13'h0521] = 0;
    assign rom[13'h0522] = 0;
    assign rom[13'h0523] = 0;
    assign rom[13'h0524] = 0;
    assign rom[13'h0525] = 0;
    assign rom[13'h0526] = 0;
    assign rom[13'h0527] = 0;
    assign rom[13'h0528] = 0;
    assign rom[13'h0529] = 0;
    assign rom[13'h052a] = 0;
    assign rom[13'h052b] = 0;
    assign rom[13'h052c] = 0;
    assign rom[13'h052d] = 0;
    assign rom[13'h052e] = 0;
    assign rom[13'h052f] = 0;
    assign rom[13'h0530] = 0;
    assign rom[13'h0531] = 0;
    assign rom[13'h0532] = 0;
    assign rom[13'h0533] = 0;
    assign rom[13'h0534] = 0;
    assign rom[13'h0535] = 0;
    assign rom[13'h0536] = 0;
    assign rom[13'h0537] = 0;
    assign rom[13'h0538] = 0;
    assign rom[13'h0539] = 0;
    assign rom[13'h053a] = 0;
    assign rom[13'h053b] = 0;
    assign rom[13'h053c] = 0;
    assign rom[13'h053d] = 0;
    assign rom[13'h053e] = 0;
    assign rom[13'h053f] = 0;
    assign rom[13'h0540] = 0;
    assign rom[13'h0541] = 0;
    assign rom[13'h0542] = 0;
    assign rom[13'h0543] = 0;
    assign rom[13'h0544] = 0;
    assign rom[13'h0545] = 0;
    assign rom[13'h0546] = 0;
    assign rom[13'h0547] = 0;
    assign rom[13'h0548] = 0;
    assign rom[13'h0549] = 0;
    assign rom[13'h054a] = 0;
    assign rom[13'h054b] = 0;
    assign rom[13'h054c] = 0;
    assign rom[13'h054d] = 0;
    assign rom[13'h054e] = 0;
    assign rom[13'h054f] = 0;
    assign rom[13'h0550] = 0;
    assign rom[13'h0551] = 0;
    assign rom[13'h0552] = 0;
    assign rom[13'h0553] = 0;
    assign rom[13'h0554] = 0;
    assign rom[13'h0555] = 0;
    assign rom[13'h0556] = 0;
    assign rom[13'h0557] = 0;
    assign rom[13'h0558] = 0;
    assign rom[13'h0559] = 0;
    assign rom[13'h055a] = 0;
    assign rom[13'h055b] = 0;
    assign rom[13'h055c] = 0;
    assign rom[13'h055d] = 0;
    assign rom[13'h055e] = 0;
    assign rom[13'h055f] = 0;
    assign rom[13'h0560] = 0;
    assign rom[13'h0561] = 0;
    assign rom[13'h0562] = 0;
    assign rom[13'h0563] = 0;
    assign rom[13'h0564] = 0;
    assign rom[13'h0565] = 0;
    assign rom[13'h0566] = 0;
    assign rom[13'h0567] = 0;
    assign rom[13'h0568] = 0;
    assign rom[13'h0569] = 0;
    assign rom[13'h056a] = 0;
    assign rom[13'h056b] = 0;
    assign rom[13'h056c] = 0;
    assign rom[13'h056d] = 0;
    assign rom[13'h056e] = 0;
    assign rom[13'h056f] = 0;
    assign rom[13'h0570] = 0;
    assign rom[13'h0571] = 0;
    assign rom[13'h0572] = 0;
    assign rom[13'h0573] = 0;
    assign rom[13'h0574] = 0;
    assign rom[13'h0575] = 0;
    assign rom[13'h0576] = 0;
    assign rom[13'h0577] = 0;
    assign rom[13'h0578] = 0;
    assign rom[13'h0579] = 0;
    assign rom[13'h057a] = 0;
    assign rom[13'h057b] = 0;
    assign rom[13'h057c] = 0;
    assign rom[13'h057d] = 0;
    assign rom[13'h057e] = 0;
    assign rom[13'h057f] = 0;
    assign rom[13'h0580] = 0;
    assign rom[13'h0581] = 0;
    assign rom[13'h0582] = 0;
    assign rom[13'h0583] = 0;
    assign rom[13'h0584] = 0;
    assign rom[13'h0585] = 0;
    assign rom[13'h0586] = 0;
    assign rom[13'h0587] = 0;
    assign rom[13'h0588] = 0;
    assign rom[13'h0589] = 0;
    assign rom[13'h058a] = 0;
    assign rom[13'h058b] = 0;
    assign rom[13'h058c] = 0;
    assign rom[13'h058d] = 0;
    assign rom[13'h058e] = 0;
    assign rom[13'h058f] = 0;
    assign rom[13'h0590] = 0;
    assign rom[13'h0591] = 0;
    assign rom[13'h0592] = 0;
    assign rom[13'h0593] = 0;
    assign rom[13'h0594] = 0;
    assign rom[13'h0595] = 0;
    assign rom[13'h0596] = 0;
    assign rom[13'h0597] = 0;
    assign rom[13'h0598] = 0;
    assign rom[13'h0599] = 0;
    assign rom[13'h059a] = 0;
    assign rom[13'h059b] = 0;
    assign rom[13'h059c] = 0;
    assign rom[13'h059d] = 0;
    assign rom[13'h059e] = 0;
    assign rom[13'h059f] = 0;
    assign rom[13'h05a0] = 0;
    assign rom[13'h05a1] = 0;
    assign rom[13'h05a2] = 0;
    assign rom[13'h05a3] = 0;
    assign rom[13'h05a4] = 0;
    assign rom[13'h05a5] = 0;
    assign rom[13'h05a6] = 0;
    assign rom[13'h05a7] = 0;
    assign rom[13'h05a8] = 0;
    assign rom[13'h05a9] = 0;
    assign rom[13'h05aa] = 0;
    assign rom[13'h05ab] = 0;
    assign rom[13'h05ac] = 0;
    assign rom[13'h05ad] = 0;
    assign rom[13'h05ae] = 0;
    assign rom[13'h05af] = 0;
    assign rom[13'h05b0] = 0;
    assign rom[13'h05b1] = 0;
    assign rom[13'h05b2] = 0;
    assign rom[13'h05b3] = 0;
    assign rom[13'h05b4] = 0;
    assign rom[13'h05b5] = 0;
    assign rom[13'h05b6] = 0;
    assign rom[13'h05b7] = 0;
    assign rom[13'h05b8] = 0;
    assign rom[13'h05b9] = 0;
    assign rom[13'h05ba] = 0;
    assign rom[13'h05bb] = 0;
    assign rom[13'h05bc] = 0;
    assign rom[13'h05bd] = 0;
    assign rom[13'h05be] = 0;
    assign rom[13'h05bf] = 0;
    assign rom[13'h05c0] = 0;
    assign rom[13'h05c1] = 0;
    assign rom[13'h05c2] = 0;
    assign rom[13'h05c3] = 0;
    assign rom[13'h05c4] = 0;
    assign rom[13'h05c5] = 0;
    assign rom[13'h05c6] = 0;
    assign rom[13'h05c7] = 0;
    assign rom[13'h05c8] = 0;
    assign rom[13'h05c9] = 0;
    assign rom[13'h05ca] = 0;
    assign rom[13'h05cb] = 0;
    assign rom[13'h05cc] = 0;
    assign rom[13'h05cd] = 0;
    assign rom[13'h05ce] = 0;
    assign rom[13'h05cf] = 0;
    assign rom[13'h05d0] = 0;
    assign rom[13'h05d1] = 0;
    assign rom[13'h05d2] = 0;
    assign rom[13'h05d3] = 0;
    assign rom[13'h05d4] = 0;
    assign rom[13'h05d5] = 0;
    assign rom[13'h05d6] = 0;
    assign rom[13'h05d7] = 0;
    assign rom[13'h05d8] = 0;
    assign rom[13'h05d9] = 0;
    assign rom[13'h05da] = 0;
    assign rom[13'h05db] = 0;
    assign rom[13'h05dc] = 0;
    assign rom[13'h05dd] = 0;
    assign rom[13'h05de] = 0;
    assign rom[13'h05df] = 0;
    assign rom[13'h05e0] = 0;
    assign rom[13'h05e1] = 0;
    assign rom[13'h05e2] = 0;
    assign rom[13'h05e3] = 0;
    assign rom[13'h05e4] = 0;
    assign rom[13'h05e5] = 0;
    assign rom[13'h05e6] = 0;
    assign rom[13'h05e7] = 0;
    assign rom[13'h05e8] = 0;
    assign rom[13'h05e9] = 0;
    assign rom[13'h05ea] = 0;
    assign rom[13'h05eb] = 0;
    assign rom[13'h05ec] = 0;
    assign rom[13'h05ed] = 0;
    assign rom[13'h05ee] = 0;
    assign rom[13'h05ef] = 0;
    assign rom[13'h05f0] = 0;
    assign rom[13'h05f1] = 0;
    assign rom[13'h05f2] = 0;
    assign rom[13'h05f3] = 0;
    assign rom[13'h05f4] = 0;
    assign rom[13'h05f5] = 0;
    assign rom[13'h05f6] = 0;
    assign rom[13'h05f7] = 0;
    assign rom[13'h05f8] = 0;
    assign rom[13'h05f9] = 0;
    assign rom[13'h05fa] = 0;
    assign rom[13'h05fb] = 0;
    assign rom[13'h05fc] = 0;
    assign rom[13'h05fd] = 0;
    assign rom[13'h05fe] = 0;
    assign rom[13'h05ff] = 0;
    assign rom[13'h0600] = 0;
    assign rom[13'h0601] = 0;
    assign rom[13'h0602] = 0;
    assign rom[13'h0603] = 0;
    assign rom[13'h0604] = 0;
    assign rom[13'h0605] = 0;
    assign rom[13'h0606] = 0;
    assign rom[13'h0607] = 0;
    assign rom[13'h0608] = 0;
    assign rom[13'h0609] = 0;
    assign rom[13'h060a] = 0;
    assign rom[13'h060b] = 0;
    assign rom[13'h060c] = 0;
    assign rom[13'h060d] = 0;
    assign rom[13'h060e] = 0;
    assign rom[13'h060f] = 0;
    assign rom[13'h0610] = 0;
    assign rom[13'h0611] = 0;
    assign rom[13'h0612] = 0;
    assign rom[13'h0613] = 0;
    assign rom[13'h0614] = 0;
    assign rom[13'h0615] = 0;
    assign rom[13'h0616] = 0;
    assign rom[13'h0617] = 0;
    assign rom[13'h0618] = 0;
    assign rom[13'h0619] = 0;
    assign rom[13'h061a] = 0;
    assign rom[13'h061b] = 0;
    assign rom[13'h061c] = 0;
    assign rom[13'h061d] = 0;
    assign rom[13'h061e] = 0;
    assign rom[13'h061f] = 0;
    assign rom[13'h0620] = 0;
    assign rom[13'h0621] = 0;
    assign rom[13'h0622] = 0;
    assign rom[13'h0623] = 0;
    assign rom[13'h0624] = 0;
    assign rom[13'h0625] = 0;
    assign rom[13'h0626] = 0;
    assign rom[13'h0627] = 0;
    assign rom[13'h0628] = 0;
    assign rom[13'h0629] = 0;
    assign rom[13'h062a] = 0;
    assign rom[13'h062b] = 0;
    assign rom[13'h062c] = 0;
    assign rom[13'h062d] = 0;
    assign rom[13'h062e] = 0;
    assign rom[13'h062f] = 0;
    assign rom[13'h0630] = 0;
    assign rom[13'h0631] = 0;
    assign rom[13'h0632] = 0;
    assign rom[13'h0633] = 0;
    assign rom[13'h0634] = 0;
    assign rom[13'h0635] = 0;
    assign rom[13'h0636] = 0;
    assign rom[13'h0637] = 0;
    assign rom[13'h0638] = 0;
    assign rom[13'h0639] = 0;
    assign rom[13'h063a] = 0;
    assign rom[13'h063b] = 0;
    assign rom[13'h063c] = 0;
    assign rom[13'h063d] = 0;
    assign rom[13'h063e] = 0;
    assign rom[13'h063f] = 0;
    assign rom[13'h0640] = 0;
    assign rom[13'h0641] = 0;
    assign rom[13'h0642] = 0;
    assign rom[13'h0643] = 0;
    assign rom[13'h0644] = 0;
    assign rom[13'h0645] = 0;
    assign rom[13'h0646] = 0;
    assign rom[13'h0647] = 0;
    assign rom[13'h0648] = 0;
    assign rom[13'h0649] = 0;
    assign rom[13'h064a] = 0;
    assign rom[13'h064b] = 0;
    assign rom[13'h064c] = 0;
    assign rom[13'h064d] = 0;
    assign rom[13'h064e] = 0;
    assign rom[13'h064f] = 0;
    assign rom[13'h0650] = 0;
    assign rom[13'h0651] = 0;
    assign rom[13'h0652] = 0;
    assign rom[13'h0653] = 0;
    assign rom[13'h0654] = 0;
    assign rom[13'h0655] = 0;
    assign rom[13'h0656] = 0;
    assign rom[13'h0657] = 0;
    assign rom[13'h0658] = 0;
    assign rom[13'h0659] = 0;
    assign rom[13'h065a] = 0;
    assign rom[13'h065b] = 0;
    assign rom[13'h065c] = 0;
    assign rom[13'h065d] = 0;
    assign rom[13'h065e] = 0;
    assign rom[13'h065f] = 0;
    assign rom[13'h0660] = 0;
    assign rom[13'h0661] = 0;
    assign rom[13'h0662] = 0;
    assign rom[13'h0663] = 0;
    assign rom[13'h0664] = 0;
    assign rom[13'h0665] = 0;
    assign rom[13'h0666] = 0;
    assign rom[13'h0667] = 0;
    assign rom[13'h0668] = 0;
    assign rom[13'h0669] = 0;
    assign rom[13'h066a] = 0;
    assign rom[13'h066b] = 0;
    assign rom[13'h066c] = 0;
    assign rom[13'h066d] = 0;
    assign rom[13'h066e] = 0;
    assign rom[13'h066f] = 0;
    assign rom[13'h0670] = 0;
    assign rom[13'h0671] = 0;
    assign rom[13'h0672] = 0;
    assign rom[13'h0673] = 0;
    assign rom[13'h0674] = 0;
    assign rom[13'h0675] = 0;
    assign rom[13'h0676] = 0;
    assign rom[13'h0677] = 0;
    assign rom[13'h0678] = 0;
    assign rom[13'h0679] = 0;
    assign rom[13'h067a] = 0;
    assign rom[13'h067b] = 0;
    assign rom[13'h067c] = 0;
    assign rom[13'h067d] = 0;
    assign rom[13'h067e] = 0;
    assign rom[13'h067f] = 0;
    assign rom[13'h0680] = 0;
    assign rom[13'h0681] = 0;
    assign rom[13'h0682] = 0;
    assign rom[13'h0683] = 0;
    assign rom[13'h0684] = 0;
    assign rom[13'h0685] = 0;
    assign rom[13'h0686] = 0;
    assign rom[13'h0687] = 0;
    assign rom[13'h0688] = 0;
    assign rom[13'h0689] = 0;
    assign rom[13'h068a] = 0;
    assign rom[13'h068b] = 0;
    assign rom[13'h068c] = 0;
    assign rom[13'h068d] = 0;
    assign rom[13'h068e] = 0;
    assign rom[13'h068f] = 0;
    assign rom[13'h0690] = 0;
    assign rom[13'h0691] = 0;
    assign rom[13'h0692] = 0;
    assign rom[13'h0693] = 0;
    assign rom[13'h0694] = 0;
    assign rom[13'h0695] = 0;
    assign rom[13'h0696] = 0;
    assign rom[13'h0697] = 0;
    assign rom[13'h0698] = 0;
    assign rom[13'h0699] = 0;
    assign rom[13'h069a] = 0;
    assign rom[13'h069b] = 0;
    assign rom[13'h069c] = 0;
    assign rom[13'h069d] = 0;
    assign rom[13'h069e] = 0;
    assign rom[13'h069f] = 0;
    assign rom[13'h06a0] = 0;
    assign rom[13'h06a1] = 0;
    assign rom[13'h06a2] = 0;
    assign rom[13'h06a3] = 0;
    assign rom[13'h06a4] = 0;
    assign rom[13'h06a5] = 0;
    assign rom[13'h06a6] = 0;
    assign rom[13'h06a7] = 0;
    assign rom[13'h06a8] = 0;
    assign rom[13'h06a9] = 0;
    assign rom[13'h06aa] = 0;
    assign rom[13'h06ab] = 0;
    assign rom[13'h06ac] = 0;
    assign rom[13'h06ad] = 0;
    assign rom[13'h06ae] = 0;
    assign rom[13'h06af] = 0;
    assign rom[13'h06b0] = 0;
    assign rom[13'h06b1] = 0;
    assign rom[13'h06b2] = 0;
    assign rom[13'h06b3] = 0;
    assign rom[13'h06b4] = 0;
    assign rom[13'h06b5] = 0;
    assign rom[13'h06b6] = 0;
    assign rom[13'h06b7] = 0;
    assign rom[13'h06b8] = 0;
    assign rom[13'h06b9] = 0;
    assign rom[13'h06ba] = 0;
    assign rom[13'h06bb] = 0;
    assign rom[13'h06bc] = 0;
    assign rom[13'h06bd] = 0;
    assign rom[13'h06be] = 0;
    assign rom[13'h06bf] = 0;
    assign rom[13'h06c0] = 0;
    assign rom[13'h06c1] = 0;
    assign rom[13'h06c2] = 0;
    assign rom[13'h06c3] = 0;
    assign rom[13'h06c4] = 0;
    assign rom[13'h06c5] = 0;
    assign rom[13'h06c6] = 0;
    assign rom[13'h06c7] = 0;
    assign rom[13'h06c8] = 0;
    assign rom[13'h06c9] = 0;
    assign rom[13'h06ca] = 0;
    assign rom[13'h06cb] = 0;
    assign rom[13'h06cc] = 0;
    assign rom[13'h06cd] = 0;
    assign rom[13'h06ce] = 0;
    assign rom[13'h06cf] = 0;
    assign rom[13'h06d0] = 0;
    assign rom[13'h06d1] = 0;
    assign rom[13'h06d2] = 0;
    assign rom[13'h06d3] = 0;
    assign rom[13'h06d4] = 0;
    assign rom[13'h06d5] = 0;
    assign rom[13'h06d6] = 0;
    assign rom[13'h06d7] = 0;
    assign rom[13'h06d8] = 0;
    assign rom[13'h06d9] = 0;
    assign rom[13'h06da] = 0;
    assign rom[13'h06db] = 0;
    assign rom[13'h06dc] = 0;
    assign rom[13'h06dd] = 0;
    assign rom[13'h06de] = 0;
    assign rom[13'h06df] = 0;
    assign rom[13'h06e0] = 0;
    assign rom[13'h06e1] = 0;
    assign rom[13'h06e2] = 0;
    assign rom[13'h06e3] = 0;
    assign rom[13'h06e4] = 0;
    assign rom[13'h06e5] = 0;
    assign rom[13'h06e6] = 0;
    assign rom[13'h06e7] = 0;
    assign rom[13'h06e8] = 0;
    assign rom[13'h06e9] = 0;
    assign rom[13'h06ea] = 0;
    assign rom[13'h06eb] = 0;
    assign rom[13'h06ec] = 0;
    assign rom[13'h06ed] = 0;
    assign rom[13'h06ee] = 0;
    assign rom[13'h06ef] = 0;
    assign rom[13'h06f0] = 0;
    assign rom[13'h06f1] = 0;
    assign rom[13'h06f2] = 0;
    assign rom[13'h06f3] = 0;
    assign rom[13'h06f4] = 0;
    assign rom[13'h06f5] = 0;
    assign rom[13'h06f6] = 0;
    assign rom[13'h06f7] = 0;
    assign rom[13'h06f8] = 0;
    assign rom[13'h06f9] = 0;
    assign rom[13'h06fa] = 0;
    assign rom[13'h06fb] = 0;
    assign rom[13'h06fc] = 0;
    assign rom[13'h06fd] = 0;
    assign rom[13'h06fe] = 0;
    assign rom[13'h06ff] = 0;
    assign rom[13'h0700] = 0;
    assign rom[13'h0701] = 0;
    assign rom[13'h0702] = 0;
    assign rom[13'h0703] = 0;
    assign rom[13'h0704] = 0;
    assign rom[13'h0705] = 0;
    assign rom[13'h0706] = 0;
    assign rom[13'h0707] = 0;
    assign rom[13'h0708] = 0;
    assign rom[13'h0709] = 0;
    assign rom[13'h070a] = 0;
    assign rom[13'h070b] = 0;
    assign rom[13'h070c] = 0;
    assign rom[13'h070d] = 0;
    assign rom[13'h070e] = 0;
    assign rom[13'h070f] = 0;
    assign rom[13'h0710] = 0;
    assign rom[13'h0711] = 0;
    assign rom[13'h0712] = 0;
    assign rom[13'h0713] = 0;
    assign rom[13'h0714] = 0;
    assign rom[13'h0715] = 0;
    assign rom[13'h0716] = 0;
    assign rom[13'h0717] = 0;
    assign rom[13'h0718] = 0;
    assign rom[13'h0719] = 0;
    assign rom[13'h071a] = 0;
    assign rom[13'h071b] = 0;
    assign rom[13'h071c] = 0;
    assign rom[13'h071d] = 0;
    assign rom[13'h071e] = 0;
    assign rom[13'h071f] = 0;
    assign rom[13'h0720] = 0;
    assign rom[13'h0721] = 0;
    assign rom[13'h0722] = 0;
    assign rom[13'h0723] = 0;
    assign rom[13'h0724] = 0;
    assign rom[13'h0725] = 0;
    assign rom[13'h0726] = 0;
    assign rom[13'h0727] = 0;
    assign rom[13'h0728] = 0;
    assign rom[13'h0729] = 0;
    assign rom[13'h072a] = 0;
    assign rom[13'h072b] = 0;
    assign rom[13'h072c] = 0;
    assign rom[13'h072d] = 0;
    assign rom[13'h072e] = 0;
    assign rom[13'h072f] = 0;
    assign rom[13'h0730] = 0;
    assign rom[13'h0731] = 0;
    assign rom[13'h0732] = 0;
    assign rom[13'h0733] = 0;
    assign rom[13'h0734] = 0;
    assign rom[13'h0735] = 0;
    assign rom[13'h0736] = 0;
    assign rom[13'h0737] = 0;
    assign rom[13'h0738] = 0;
    assign rom[13'h0739] = 0;
    assign rom[13'h073a] = 0;
    assign rom[13'h073b] = 0;
    assign rom[13'h073c] = 0;
    assign rom[13'h073d] = 0;
    assign rom[13'h073e] = 0;
    assign rom[13'h073f] = 0;
    assign rom[13'h0740] = 0;
    assign rom[13'h0741] = 0;
    assign rom[13'h0742] = 0;
    assign rom[13'h0743] = 0;
    assign rom[13'h0744] = 0;
    assign rom[13'h0745] = 0;
    assign rom[13'h0746] = 0;
    assign rom[13'h0747] = 0;
    assign rom[13'h0748] = 0;
    assign rom[13'h0749] = 0;
    assign rom[13'h074a] = 0;
    assign rom[13'h074b] = 0;
    assign rom[13'h074c] = 0;
    assign rom[13'h074d] = 0;
    assign rom[13'h074e] = 0;
    assign rom[13'h074f] = 0;
    assign rom[13'h0750] = 0;
    assign rom[13'h0751] = 0;
    assign rom[13'h0752] = 0;
    assign rom[13'h0753] = 0;
    assign rom[13'h0754] = 0;
    assign rom[13'h0755] = 0;
    assign rom[13'h0756] = 0;
    assign rom[13'h0757] = 0;
    assign rom[13'h0758] = 0;
    assign rom[13'h0759] = 0;
    assign rom[13'h075a] = 0;
    assign rom[13'h075b] = 0;
    assign rom[13'h075c] = 0;
    assign rom[13'h075d] = 0;
    assign rom[13'h075e] = 0;
    assign rom[13'h075f] = 0;
    assign rom[13'h0760] = 0;
    assign rom[13'h0761] = 0;
    assign rom[13'h0762] = 0;
    assign rom[13'h0763] = 0;
    assign rom[13'h0764] = 0;
    assign rom[13'h0765] = 0;
    assign rom[13'h0766] = 0;
    assign rom[13'h0767] = 0;
    assign rom[13'h0768] = 0;
    assign rom[13'h0769] = 0;
    assign rom[13'h076a] = 0;
    assign rom[13'h076b] = 0;
    assign rom[13'h076c] = 0;
    assign rom[13'h076d] = 0;
    assign rom[13'h076e] = 0;
    assign rom[13'h076f] = 0;
    assign rom[13'h0770] = 0;
    assign rom[13'h0771] = 0;
    assign rom[13'h0772] = 0;
    assign rom[13'h0773] = 0;
    assign rom[13'h0774] = 0;
    assign rom[13'h0775] = 0;
    assign rom[13'h0776] = 0;
    assign rom[13'h0777] = 0;
    assign rom[13'h0778] = 0;
    assign rom[13'h0779] = 0;
    assign rom[13'h077a] = 0;
    assign rom[13'h077b] = 0;
    assign rom[13'h077c] = 0;
    assign rom[13'h077d] = 0;
    assign rom[13'h077e] = 0;
    assign rom[13'h077f] = 0;
    assign rom[13'h0780] = 0;
    assign rom[13'h0781] = 0;
    assign rom[13'h0782] = 0;
    assign rom[13'h0783] = 0;
    assign rom[13'h0784] = 0;
    assign rom[13'h0785] = 0;
    assign rom[13'h0786] = 0;
    assign rom[13'h0787] = 0;
    assign rom[13'h0788] = 0;
    assign rom[13'h0789] = 0;
    assign rom[13'h078a] = 0;
    assign rom[13'h078b] = 0;
    assign rom[13'h078c] = 0;
    assign rom[13'h078d] = 0;
    assign rom[13'h078e] = 0;
    assign rom[13'h078f] = 0;
    assign rom[13'h0790] = 0;
    assign rom[13'h0791] = 0;
    assign rom[13'h0792] = 0;
    assign rom[13'h0793] = 0;
    assign rom[13'h0794] = 0;
    assign rom[13'h0795] = 0;
    assign rom[13'h0796] = 0;
    assign rom[13'h0797] = 0;
    assign rom[13'h0798] = 0;
    assign rom[13'h0799] = 0;
    assign rom[13'h079a] = 0;
    assign rom[13'h079b] = 0;
    assign rom[13'h079c] = 0;
    assign rom[13'h079d] = 0;
    assign rom[13'h079e] = 0;
    assign rom[13'h079f] = 0;
    assign rom[13'h07a0] = 0;
    assign rom[13'h07a1] = 0;
    assign rom[13'h07a2] = 0;
    assign rom[13'h07a3] = 0;
    assign rom[13'h07a4] = 0;
    assign rom[13'h07a5] = 0;
    assign rom[13'h07a6] = 0;
    assign rom[13'h07a7] = 0;
    assign rom[13'h07a8] = 0;
    assign rom[13'h07a9] = 0;
    assign rom[13'h07aa] = 0;
    assign rom[13'h07ab] = 0;
    assign rom[13'h07ac] = 0;
    assign rom[13'h07ad] = 0;
    assign rom[13'h07ae] = 0;
    assign rom[13'h07af] = 0;
    assign rom[13'h07b0] = 0;
    assign rom[13'h07b1] = 0;
    assign rom[13'h07b2] = 0;
    assign rom[13'h07b3] = 0;
    assign rom[13'h07b4] = 0;
    assign rom[13'h07b5] = 0;
    assign rom[13'h07b6] = 0;
    assign rom[13'h07b7] = 0;
    assign rom[13'h07b8] = 0;
    assign rom[13'h07b9] = 0;
    assign rom[13'h07ba] = 0;
    assign rom[13'h07bb] = 0;
    assign rom[13'h07bc] = 0;
    assign rom[13'h07bd] = 0;
    assign rom[13'h07be] = 0;
    assign rom[13'h07bf] = 0;
    assign rom[13'h07c0] = 0;
    assign rom[13'h07c1] = 0;
    assign rom[13'h07c2] = 0;
    assign rom[13'h07c3] = 0;
    assign rom[13'h07c4] = 0;
    assign rom[13'h07c5] = 0;
    assign rom[13'h07c6] = 0;
    assign rom[13'h07c7] = 0;
    assign rom[13'h07c8] = 0;
    assign rom[13'h07c9] = 0;
    assign rom[13'h07ca] = 0;
    assign rom[13'h07cb] = 0;
    assign rom[13'h07cc] = 0;
    assign rom[13'h07cd] = 0;
    assign rom[13'h07ce] = 0;
    assign rom[13'h07cf] = 0;
    assign rom[13'h07d0] = 0;
    assign rom[13'h07d1] = 0;
    assign rom[13'h07d2] = 0;
    assign rom[13'h07d3] = 0;
    assign rom[13'h07d4] = 0;
    assign rom[13'h07d5] = 0;
    assign rom[13'h07d6] = 0;
    assign rom[13'h07d7] = 0;
    assign rom[13'h07d8] = 0;
    assign rom[13'h07d9] = 0;
    assign rom[13'h07da] = 0;
    assign rom[13'h07db] = 0;
    assign rom[13'h07dc] = 0;
    assign rom[13'h07dd] = 0;
    assign rom[13'h07de] = 0;
    assign rom[13'h07df] = 0;
    assign rom[13'h07e0] = 0;
    assign rom[13'h07e1] = 0;
    assign rom[13'h07e2] = 0;
    assign rom[13'h07e3] = 0;
    assign rom[13'h07e4] = 0;
    assign rom[13'h07e5] = 0;
    assign rom[13'h07e6] = 0;
    assign rom[13'h07e7] = 0;
    assign rom[13'h07e8] = 0;
    assign rom[13'h07e9] = 0;
    assign rom[13'h07ea] = 0;
    assign rom[13'h07eb] = 0;
    assign rom[13'h07ec] = 0;
    assign rom[13'h07ed] = 0;
    assign rom[13'h07ee] = 0;
    assign rom[13'h07ef] = 0;
    assign rom[13'h07f0] = 0;
    assign rom[13'h07f1] = 0;
    assign rom[13'h07f2] = 0;
    assign rom[13'h07f3] = 0;
    assign rom[13'h07f4] = 0;
    assign rom[13'h07f5] = 0;
    assign rom[13'h07f6] = 0;
    assign rom[13'h07f7] = 0;
    assign rom[13'h07f8] = 0;
    assign rom[13'h07f9] = 0;
    assign rom[13'h07fa] = 0;
    assign rom[13'h07fb] = 0;
    assign rom[13'h07fc] = 0;
    assign rom[13'h07fd] = 0;
    assign rom[13'h07fe] = 0;
    assign rom[13'h07ff] = 0;
    assign rom[13'h0800] = 0;
    assign rom[13'h0801] = 0;
    assign rom[13'h0802] = 0;
    assign rom[13'h0803] = 0;
    assign rom[13'h0804] = 0;
    assign rom[13'h0805] = 0;
    assign rom[13'h0806] = 0;
    assign rom[13'h0807] = 0;
    assign rom[13'h0808] = 0;
    assign rom[13'h0809] = 0;
    assign rom[13'h080a] = 0;
    assign rom[13'h080b] = 0;
    assign rom[13'h080c] = 0;
    assign rom[13'h080d] = 0;
    assign rom[13'h080e] = 0;
    assign rom[13'h080f] = 0;
    assign rom[13'h0810] = 0;
    assign rom[13'h0811] = 0;
    assign rom[13'h0812] = 0;
    assign rom[13'h0813] = 0;
    assign rom[13'h0814] = 0;
    assign rom[13'h0815] = 0;
    assign rom[13'h0816] = 0;
    assign rom[13'h0817] = 0;
    assign rom[13'h0818] = 0;
    assign rom[13'h0819] = 0;
    assign rom[13'h081a] = 0;
    assign rom[13'h081b] = 0;
    assign rom[13'h081c] = 0;
    assign rom[13'h081d] = 0;
    assign rom[13'h081e] = 0;
    assign rom[13'h081f] = 0;
    assign rom[13'h0820] = 0;
    assign rom[13'h0821] = 0;
    assign rom[13'h0822] = 0;
    assign rom[13'h0823] = 0;
    assign rom[13'h0824] = 0;
    assign rom[13'h0825] = 0;
    assign rom[13'h0826] = 0;
    assign rom[13'h0827] = 0;
    assign rom[13'h0828] = 0;
    assign rom[13'h0829] = 0;
    assign rom[13'h082a] = 0;
    assign rom[13'h082b] = 0;
    assign rom[13'h082c] = 0;
    assign rom[13'h082d] = 0;
    assign rom[13'h082e] = 0;
    assign rom[13'h082f] = 0;
    assign rom[13'h0830] = 0;
    assign rom[13'h0831] = 0;
    assign rom[13'h0832] = 0;
    assign rom[13'h0833] = 0;
    assign rom[13'h0834] = 0;
    assign rom[13'h0835] = 0;
    assign rom[13'h0836] = 0;
    assign rom[13'h0837] = 0;
    assign rom[13'h0838] = 0;
    assign rom[13'h0839] = 0;
    assign rom[13'h083a] = 0;
    assign rom[13'h083b] = 0;
    assign rom[13'h083c] = 0;
    assign rom[13'h083d] = 0;
    assign rom[13'h083e] = 0;
    assign rom[13'h083f] = 0;
    assign rom[13'h0840] = 0;
    assign rom[13'h0841] = 0;
    assign rom[13'h0842] = 0;
    assign rom[13'h0843] = 1;
    assign rom[13'h0844] = 1;
    assign rom[13'h0845] = 0;
    assign rom[13'h0846] = 0;
    assign rom[13'h0847] = 0;
    assign rom[13'h0848] = 0;
    assign rom[13'h0849] = 0;
    assign rom[13'h084a] = 0;
    assign rom[13'h084b] = 1;
    assign rom[13'h084c] = 1;
    assign rom[13'h084d] = 0;
    assign rom[13'h084e] = 0;
    assign rom[13'h084f] = 0;
    assign rom[13'h0850] = 0;
    assign rom[13'h0851] = 0;
    assign rom[13'h0852] = 0;
    assign rom[13'h0853] = 1;
    assign rom[13'h0854] = 1;
    assign rom[13'h0855] = 0;
    assign rom[13'h0856] = 0;
    assign rom[13'h0857] = 0;
    assign rom[13'h0858] = 0;
    assign rom[13'h0859] = 0;
    assign rom[13'h085a] = 0;
    assign rom[13'h085b] = 1;
    assign rom[13'h085c] = 1;
    assign rom[13'h085d] = 0;
    assign rom[13'h085e] = 0;
    assign rom[13'h085f] = 0;
    assign rom[13'h0860] = 0;
    assign rom[13'h0861] = 0;
    assign rom[13'h0862] = 0;
    assign rom[13'h0863] = 0;
    assign rom[13'h0864] = 0;
    assign rom[13'h0865] = 0;
    assign rom[13'h0866] = 0;
    assign rom[13'h0867] = 0;
    assign rom[13'h0868] = 0;
    assign rom[13'h0869] = 0;
    assign rom[13'h086a] = 0;
    assign rom[13'h086b] = 1;
    assign rom[13'h086c] = 1;
    assign rom[13'h086d] = 0;
    assign rom[13'h086e] = 0;
    assign rom[13'h086f] = 0;
    assign rom[13'h0870] = 0;
    assign rom[13'h0871] = 0;
    assign rom[13'h0872] = 0;
    assign rom[13'h0873] = 1;
    assign rom[13'h0874] = 1;
    assign rom[13'h0875] = 0;
    assign rom[13'h0876] = 0;
    assign rom[13'h0877] = 0;
    assign rom[13'h0878] = 0;
    assign rom[13'h0879] = 0;
    assign rom[13'h087a] = 0;
    assign rom[13'h087b] = 0;
    assign rom[13'h087c] = 0;
    assign rom[13'h087d] = 0;
    assign rom[13'h087e] = 0;
    assign rom[13'h087f] = 0;
    assign rom[13'h0880] = 0;
    assign rom[13'h0881] = 1;
    assign rom[13'h0882] = 1;
    assign rom[13'h0883] = 0;
    assign rom[13'h0884] = 1;
    assign rom[13'h0885] = 1;
    assign rom[13'h0886] = 0;
    assign rom[13'h0887] = 0;
    assign rom[13'h0888] = 0;
    assign rom[13'h0889] = 1;
    assign rom[13'h088a] = 1;
    assign rom[13'h088b] = 0;
    assign rom[13'h088c] = 1;
    assign rom[13'h088d] = 1;
    assign rom[13'h088e] = 0;
    assign rom[13'h088f] = 0;
    assign rom[13'h0890] = 0;
    assign rom[13'h0891] = 1;
    assign rom[13'h0892] = 0;
    assign rom[13'h0893] = 0;
    assign rom[13'h0894] = 1;
    assign rom[13'h0895] = 0;
    assign rom[13'h0896] = 0;
    assign rom[13'h0897] = 0;
    assign rom[13'h0898] = 0;
    assign rom[13'h0899] = 0;
    assign rom[13'h089a] = 0;
    assign rom[13'h089b] = 0;
    assign rom[13'h089c] = 0;
    assign rom[13'h089d] = 0;
    assign rom[13'h089e] = 0;
    assign rom[13'h089f] = 0;
    assign rom[13'h08a0] = 0;
    assign rom[13'h08a1] = 0;
    assign rom[13'h08a2] = 0;
    assign rom[13'h08a3] = 0;
    assign rom[13'h08a4] = 0;
    assign rom[13'h08a5] = 0;
    assign rom[13'h08a6] = 0;
    assign rom[13'h08a7] = 0;
    assign rom[13'h08a8] = 0;
    assign rom[13'h08a9] = 0;
    assign rom[13'h08aa] = 0;
    assign rom[13'h08ab] = 0;
    assign rom[13'h08ac] = 0;
    assign rom[13'h08ad] = 0;
    assign rom[13'h08ae] = 0;
    assign rom[13'h08af] = 0;
    assign rom[13'h08b0] = 0;
    assign rom[13'h08b1] = 0;
    assign rom[13'h08b2] = 0;
    assign rom[13'h08b3] = 0;
    assign rom[13'h08b4] = 0;
    assign rom[13'h08b5] = 0;
    assign rom[13'h08b6] = 0;
    assign rom[13'h08b7] = 0;
    assign rom[13'h08b8] = 0;
    assign rom[13'h08b9] = 0;
    assign rom[13'h08ba] = 0;
    assign rom[13'h08bb] = 0;
    assign rom[13'h08bc] = 0;
    assign rom[13'h08bd] = 0;
    assign rom[13'h08be] = 0;
    assign rom[13'h08bf] = 0;
    assign rom[13'h08c0] = 0;
    assign rom[13'h08c1] = 1;
    assign rom[13'h08c2] = 1;
    assign rom[13'h08c3] = 0;
    assign rom[13'h08c4] = 1;
    assign rom[13'h08c5] = 1;
    assign rom[13'h08c6] = 0;
    assign rom[13'h08c7] = 0;
    assign rom[13'h08c8] = 0;
    assign rom[13'h08c9] = 1;
    assign rom[13'h08ca] = 1;
    assign rom[13'h08cb] = 0;
    assign rom[13'h08cc] = 1;
    assign rom[13'h08cd] = 1;
    assign rom[13'h08ce] = 0;
    assign rom[13'h08cf] = 0;
    assign rom[13'h08d0] = 1;
    assign rom[13'h08d1] = 1;
    assign rom[13'h08d2] = 1;
    assign rom[13'h08d3] = 1;
    assign rom[13'h08d4] = 1;
    assign rom[13'h08d5] = 1;
    assign rom[13'h08d6] = 1;
    assign rom[13'h08d7] = 0;
    assign rom[13'h08d8] = 0;
    assign rom[13'h08d9] = 1;
    assign rom[13'h08da] = 1;
    assign rom[13'h08db] = 0;
    assign rom[13'h08dc] = 1;
    assign rom[13'h08dd] = 1;
    assign rom[13'h08de] = 0;
    assign rom[13'h08df] = 0;
    assign rom[13'h08e0] = 1;
    assign rom[13'h08e1] = 1;
    assign rom[13'h08e2] = 1;
    assign rom[13'h08e3] = 1;
    assign rom[13'h08e4] = 1;
    assign rom[13'h08e5] = 1;
    assign rom[13'h08e6] = 1;
    assign rom[13'h08e7] = 0;
    assign rom[13'h08e8] = 0;
    assign rom[13'h08e9] = 1;
    assign rom[13'h08ea] = 1;
    assign rom[13'h08eb] = 0;
    assign rom[13'h08ec] = 1;
    assign rom[13'h08ed] = 1;
    assign rom[13'h08ee] = 0;
    assign rom[13'h08ef] = 0;
    assign rom[13'h08f0] = 0;
    assign rom[13'h08f1] = 1;
    assign rom[13'h08f2] = 1;
    assign rom[13'h08f3] = 0;
    assign rom[13'h08f4] = 1;
    assign rom[13'h08f5] = 1;
    assign rom[13'h08f6] = 0;
    assign rom[13'h08f7] = 0;
    assign rom[13'h08f8] = 0;
    assign rom[13'h08f9] = 0;
    assign rom[13'h08fa] = 0;
    assign rom[13'h08fb] = 0;
    assign rom[13'h08fc] = 0;
    assign rom[13'h08fd] = 0;
    assign rom[13'h08fe] = 0;
    assign rom[13'h08ff] = 0;
    assign rom[13'h0900] = 0;
    assign rom[13'h0901] = 0;
    assign rom[13'h0902] = 0;
    assign rom[13'h0903] = 1;
    assign rom[13'h0904] = 1;
    assign rom[13'h0905] = 0;
    assign rom[13'h0906] = 0;
    assign rom[13'h0907] = 0;
    assign rom[13'h0908] = 0;
    assign rom[13'h0909] = 1;
    assign rom[13'h090a] = 1;
    assign rom[13'h090b] = 1;
    assign rom[13'h090c] = 1;
    assign rom[13'h090d] = 1;
    assign rom[13'h090e] = 1;
    assign rom[13'h090f] = 0;
    assign rom[13'h0910] = 1;
    assign rom[13'h0911] = 1;
    assign rom[13'h0912] = 0;
    assign rom[13'h0913] = 1;
    assign rom[13'h0914] = 1;
    assign rom[13'h0915] = 0;
    assign rom[13'h0916] = 0;
    assign rom[13'h0917] = 0;
    assign rom[13'h0918] = 0;
    assign rom[13'h0919] = 1;
    assign rom[13'h091a] = 1;
    assign rom[13'h091b] = 1;
    assign rom[13'h091c] = 1;
    assign rom[13'h091d] = 1;
    assign rom[13'h091e] = 1;
    assign rom[13'h091f] = 0;
    assign rom[13'h0920] = 0;
    assign rom[13'h0921] = 0;
    assign rom[13'h0922] = 0;
    assign rom[13'h0923] = 1;
    assign rom[13'h0924] = 1;
    assign rom[13'h0925] = 0;
    assign rom[13'h0926] = 1;
    assign rom[13'h0927] = 1;
    assign rom[13'h0928] = 0;
    assign rom[13'h0929] = 1;
    assign rom[13'h092a] = 1;
    assign rom[13'h092b] = 1;
    assign rom[13'h092c] = 1;
    assign rom[13'h092d] = 1;
    assign rom[13'h092e] = 1;
    assign rom[13'h092f] = 0;
    assign rom[13'h0930] = 0;
    assign rom[13'h0931] = 0;
    assign rom[13'h0932] = 0;
    assign rom[13'h0933] = 1;
    assign rom[13'h0934] = 1;
    assign rom[13'h0935] = 0;
    assign rom[13'h0936] = 0;
    assign rom[13'h0937] = 0;
    assign rom[13'h0938] = 0;
    assign rom[13'h0939] = 0;
    assign rom[13'h093a] = 0;
    assign rom[13'h093b] = 0;
    assign rom[13'h093c] = 0;
    assign rom[13'h093d] = 0;
    assign rom[13'h093e] = 0;
    assign rom[13'h093f] = 0;
    assign rom[13'h0940] = 0;
    assign rom[13'h0941] = 1;
    assign rom[13'h0942] = 1;
    assign rom[13'h0943] = 0;
    assign rom[13'h0944] = 0;
    assign rom[13'h0945] = 0;
    assign rom[13'h0946] = 1;
    assign rom[13'h0947] = 0;
    assign rom[13'h0948] = 0;
    assign rom[13'h0949] = 1;
    assign rom[13'h094a] = 1;
    assign rom[13'h094b] = 0;
    assign rom[13'h094c] = 0;
    assign rom[13'h094d] = 1;
    assign rom[13'h094e] = 1;
    assign rom[13'h094f] = 0;
    assign rom[13'h0950] = 0;
    assign rom[13'h0951] = 0;
    assign rom[13'h0952] = 0;
    assign rom[13'h0953] = 0;
    assign rom[13'h0954] = 1;
    assign rom[13'h0955] = 1;
    assign rom[13'h0956] = 0;
    assign rom[13'h0957] = 0;
    assign rom[13'h0958] = 0;
    assign rom[13'h0959] = 0;
    assign rom[13'h095a] = 0;
    assign rom[13'h095b] = 1;
    assign rom[13'h095c] = 1;
    assign rom[13'h095d] = 0;
    assign rom[13'h095e] = 0;
    assign rom[13'h095f] = 0;
    assign rom[13'h0960] = 0;
    assign rom[13'h0961] = 0;
    assign rom[13'h0962] = 1;
    assign rom[13'h0963] = 1;
    assign rom[13'h0964] = 0;
    assign rom[13'h0965] = 0;
    assign rom[13'h0966] = 0;
    assign rom[13'h0967] = 0;
    assign rom[13'h0968] = 0;
    assign rom[13'h0969] = 1;
    assign rom[13'h096a] = 1;
    assign rom[13'h096b] = 0;
    assign rom[13'h096c] = 0;
    assign rom[13'h096d] = 1;
    assign rom[13'h096e] = 1;
    assign rom[13'h096f] = 0;
    assign rom[13'h0970] = 0;
    assign rom[13'h0971] = 1;
    assign rom[13'h0972] = 0;
    assign rom[13'h0973] = 0;
    assign rom[13'h0974] = 0;
    assign rom[13'h0975] = 1;
    assign rom[13'h0976] = 1;
    assign rom[13'h0977] = 0;
    assign rom[13'h0978] = 0;
    assign rom[13'h0979] = 0;
    assign rom[13'h097a] = 0;
    assign rom[13'h097b] = 0;
    assign rom[13'h097c] = 0;
    assign rom[13'h097d] = 0;
    assign rom[13'h097e] = 0;
    assign rom[13'h097f] = 0;
    assign rom[13'h0980] = 0;
    assign rom[13'h0981] = 0;
    assign rom[13'h0982] = 1;
    assign rom[13'h0983] = 1;
    assign rom[13'h0984] = 1;
    assign rom[13'h0985] = 0;
    assign rom[13'h0986] = 0;
    assign rom[13'h0987] = 0;
    assign rom[13'h0988] = 0;
    assign rom[13'h0989] = 1;
    assign rom[13'h098a] = 1;
    assign rom[13'h098b] = 0;
    assign rom[13'h098c] = 1;
    assign rom[13'h098d] = 1;
    assign rom[13'h098e] = 0;
    assign rom[13'h098f] = 0;
    assign rom[13'h0990] = 0;
    assign rom[13'h0991] = 1;
    assign rom[13'h0992] = 1;
    assign rom[13'h0993] = 0;
    assign rom[13'h0994] = 1;
    assign rom[13'h0995] = 0;
    assign rom[13'h0996] = 0;
    assign rom[13'h0997] = 0;
    assign rom[13'h0998] = 0;
    assign rom[13'h0999] = 1;
    assign rom[13'h099a] = 1;
    assign rom[13'h099b] = 1;
    assign rom[13'h099c] = 0;
    assign rom[13'h099d] = 1;
    assign rom[13'h099e] = 1;
    assign rom[13'h099f] = 0;
    assign rom[13'h09a0] = 1;
    assign rom[13'h09a1] = 1;
    assign rom[13'h09a2] = 0;
    assign rom[13'h09a3] = 1;
    assign rom[13'h09a4] = 1;
    assign rom[13'h09a5] = 1;
    assign rom[13'h09a6] = 0;
    assign rom[13'h09a7] = 0;
    assign rom[13'h09a8] = 1;
    assign rom[13'h09a9] = 1;
    assign rom[13'h09aa] = 0;
    assign rom[13'h09ab] = 0;
    assign rom[13'h09ac] = 1;
    assign rom[13'h09ad] = 1;
    assign rom[13'h09ae] = 0;
    assign rom[13'h09af] = 0;
    assign rom[13'h09b0] = 0;
    assign rom[13'h09b1] = 1;
    assign rom[13'h09b2] = 1;
    assign rom[13'h09b3] = 1;
    assign rom[13'h09b4] = 0;
    assign rom[13'h09b5] = 1;
    assign rom[13'h09b6] = 1;
    assign rom[13'h09b7] = 0;
    assign rom[13'h09b8] = 0;
    assign rom[13'h09b9] = 0;
    assign rom[13'h09ba] = 0;
    assign rom[13'h09bb] = 0;
    assign rom[13'h09bc] = 0;
    assign rom[13'h09bd] = 0;
    assign rom[13'h09be] = 0;
    assign rom[13'h09bf] = 0;
    assign rom[13'h09c0] = 0;
    assign rom[13'h09c1] = 0;
    assign rom[13'h09c2] = 0;
    assign rom[13'h09c3] = 1;
    assign rom[13'h09c4] = 1;
    assign rom[13'h09c5] = 0;
    assign rom[13'h09c6] = 0;
    assign rom[13'h09c7] = 0;
    assign rom[13'h09c8] = 0;
    assign rom[13'h09c9] = 0;
    assign rom[13'h09ca] = 0;
    assign rom[13'h09cb] = 1;
    assign rom[13'h09cc] = 1;
    assign rom[13'h09cd] = 0;
    assign rom[13'h09ce] = 0;
    assign rom[13'h09cf] = 0;
    assign rom[13'h09d0] = 0;
    assign rom[13'h09d1] = 0;
    assign rom[13'h09d2] = 1;
    assign rom[13'h09d3] = 1;
    assign rom[13'h09d4] = 0;
    assign rom[13'h09d5] = 0;
    assign rom[13'h09d6] = 0;
    assign rom[13'h09d7] = 0;
    assign rom[13'h09d8] = 0;
    assign rom[13'h09d9] = 0;
    assign rom[13'h09da] = 0;
    assign rom[13'h09db] = 0;
    assign rom[13'h09dc] = 0;
    assign rom[13'h09dd] = 0;
    assign rom[13'h09de] = 0;
    assign rom[13'h09df] = 0;
    assign rom[13'h09e0] = 0;
    assign rom[13'h09e1] = 0;
    assign rom[13'h09e2] = 0;
    assign rom[13'h09e3] = 0;
    assign rom[13'h09e4] = 0;
    assign rom[13'h09e5] = 0;
    assign rom[13'h09e6] = 0;
    assign rom[13'h09e7] = 0;
    assign rom[13'h09e8] = 0;
    assign rom[13'h09e9] = 0;
    assign rom[13'h09ea] = 0;
    assign rom[13'h09eb] = 0;
    assign rom[13'h09ec] = 0;
    assign rom[13'h09ed] = 0;
    assign rom[13'h09ee] = 0;
    assign rom[13'h09ef] = 0;
    assign rom[13'h09f0] = 0;
    assign rom[13'h09f1] = 0;
    assign rom[13'h09f2] = 0;
    assign rom[13'h09f3] = 0;
    assign rom[13'h09f4] = 0;
    assign rom[13'h09f5] = 0;
    assign rom[13'h09f6] = 0;
    assign rom[13'h09f7] = 0;
    assign rom[13'h09f8] = 0;
    assign rom[13'h09f9] = 0;
    assign rom[13'h09fa] = 0;
    assign rom[13'h09fb] = 0;
    assign rom[13'h09fc] = 0;
    assign rom[13'h09fd] = 0;
    assign rom[13'h09fe] = 0;
    assign rom[13'h09ff] = 0;
    assign rom[13'h0a00] = 0;
    assign rom[13'h0a01] = 0;
    assign rom[13'h0a02] = 0;
    assign rom[13'h0a03] = 0;
    assign rom[13'h0a04] = 1;
    assign rom[13'h0a05] = 1;
    assign rom[13'h0a06] = 0;
    assign rom[13'h0a07] = 0;
    assign rom[13'h0a08] = 0;
    assign rom[13'h0a09] = 0;
    assign rom[13'h0a0a] = 0;
    assign rom[13'h0a0b] = 1;
    assign rom[13'h0a0c] = 1;
    assign rom[13'h0a0d] = 0;
    assign rom[13'h0a0e] = 0;
    assign rom[13'h0a0f] = 0;
    assign rom[13'h0a10] = 0;
    assign rom[13'h0a11] = 0;
    assign rom[13'h0a12] = 1;
    assign rom[13'h0a13] = 1;
    assign rom[13'h0a14] = 0;
    assign rom[13'h0a15] = 0;
    assign rom[13'h0a16] = 0;
    assign rom[13'h0a17] = 0;
    assign rom[13'h0a18] = 0;
    assign rom[13'h0a19] = 0;
    assign rom[13'h0a1a] = 1;
    assign rom[13'h0a1b] = 1;
    assign rom[13'h0a1c] = 0;
    assign rom[13'h0a1d] = 0;
    assign rom[13'h0a1e] = 0;
    assign rom[13'h0a1f] = 0;
    assign rom[13'h0a20] = 0;
    assign rom[13'h0a21] = 0;
    assign rom[13'h0a22] = 1;
    assign rom[13'h0a23] = 1;
    assign rom[13'h0a24] = 0;
    assign rom[13'h0a25] = 0;
    assign rom[13'h0a26] = 0;
    assign rom[13'h0a27] = 0;
    assign rom[13'h0a28] = 0;
    assign rom[13'h0a29] = 0;
    assign rom[13'h0a2a] = 0;
    assign rom[13'h0a2b] = 1;
    assign rom[13'h0a2c] = 1;
    assign rom[13'h0a2d] = 0;
    assign rom[13'h0a2e] = 0;
    assign rom[13'h0a2f] = 0;
    assign rom[13'h0a30] = 0;
    assign rom[13'h0a31] = 0;
    assign rom[13'h0a32] = 0;
    assign rom[13'h0a33] = 0;
    assign rom[13'h0a34] = 1;
    assign rom[13'h0a35] = 1;
    assign rom[13'h0a36] = 0;
    assign rom[13'h0a37] = 0;
    assign rom[13'h0a38] = 0;
    assign rom[13'h0a39] = 0;
    assign rom[13'h0a3a] = 0;
    assign rom[13'h0a3b] = 0;
    assign rom[13'h0a3c] = 0;
    assign rom[13'h0a3d] = 0;
    assign rom[13'h0a3e] = 0;
    assign rom[13'h0a3f] = 0;
    assign rom[13'h0a40] = 0;
    assign rom[13'h0a41] = 0;
    assign rom[13'h0a42] = 1;
    assign rom[13'h0a43] = 1;
    assign rom[13'h0a44] = 0;
    assign rom[13'h0a45] = 0;
    assign rom[13'h0a46] = 0;
    assign rom[13'h0a47] = 0;
    assign rom[13'h0a48] = 0;
    assign rom[13'h0a49] = 0;
    assign rom[13'h0a4a] = 0;
    assign rom[13'h0a4b] = 1;
    assign rom[13'h0a4c] = 1;
    assign rom[13'h0a4d] = 0;
    assign rom[13'h0a4e] = 0;
    assign rom[13'h0a4f] = 0;
    assign rom[13'h0a50] = 0;
    assign rom[13'h0a51] = 0;
    assign rom[13'h0a52] = 0;
    assign rom[13'h0a53] = 0;
    assign rom[13'h0a54] = 1;
    assign rom[13'h0a55] = 1;
    assign rom[13'h0a56] = 0;
    assign rom[13'h0a57] = 0;
    assign rom[13'h0a58] = 0;
    assign rom[13'h0a59] = 0;
    assign rom[13'h0a5a] = 0;
    assign rom[13'h0a5b] = 0;
    assign rom[13'h0a5c] = 1;
    assign rom[13'h0a5d] = 1;
    assign rom[13'h0a5e] = 0;
    assign rom[13'h0a5f] = 0;
    assign rom[13'h0a60] = 0;
    assign rom[13'h0a61] = 0;
    assign rom[13'h0a62] = 0;
    assign rom[13'h0a63] = 0;
    assign rom[13'h0a64] = 1;
    assign rom[13'h0a65] = 1;
    assign rom[13'h0a66] = 0;
    assign rom[13'h0a67] = 0;
    assign rom[13'h0a68] = 0;
    assign rom[13'h0a69] = 0;
    assign rom[13'h0a6a] = 0;
    assign rom[13'h0a6b] = 1;
    assign rom[13'h0a6c] = 1;
    assign rom[13'h0a6d] = 0;
    assign rom[13'h0a6e] = 0;
    assign rom[13'h0a6f] = 0;
    assign rom[13'h0a70] = 0;
    assign rom[13'h0a71] = 0;
    assign rom[13'h0a72] = 1;
    assign rom[13'h0a73] = 1;
    assign rom[13'h0a74] = 0;
    assign rom[13'h0a75] = 0;
    assign rom[13'h0a76] = 0;
    assign rom[13'h0a77] = 0;
    assign rom[13'h0a78] = 0;
    assign rom[13'h0a79] = 0;
    assign rom[13'h0a7a] = 0;
    assign rom[13'h0a7b] = 0;
    assign rom[13'h0a7c] = 0;
    assign rom[13'h0a7d] = 0;
    assign rom[13'h0a7e] = 0;
    assign rom[13'h0a7f] = 0;
    assign rom[13'h0a80] = 0;
    assign rom[13'h0a81] = 0;
    assign rom[13'h0a82] = 0;
    assign rom[13'h0a83] = 0;
    assign rom[13'h0a84] = 0;
    assign rom[13'h0a85] = 0;
    assign rom[13'h0a86] = 0;
    assign rom[13'h0a87] = 0;
    assign rom[13'h0a88] = 0;
    assign rom[13'h0a89] = 1;
    assign rom[13'h0a8a] = 1;
    assign rom[13'h0a8b] = 0;
    assign rom[13'h0a8c] = 1;
    assign rom[13'h0a8d] = 1;
    assign rom[13'h0a8e] = 0;
    assign rom[13'h0a8f] = 0;
    assign rom[13'h0a90] = 0;
    assign rom[13'h0a91] = 0;
    assign rom[13'h0a92] = 1;
    assign rom[13'h0a93] = 1;
    assign rom[13'h0a94] = 1;
    assign rom[13'h0a95] = 0;
    assign rom[13'h0a96] = 0;
    assign rom[13'h0a97] = 0;
    assign rom[13'h0a98] = 1;
    assign rom[13'h0a99] = 1;
    assign rom[13'h0a9a] = 1;
    assign rom[13'h0a9b] = 1;
    assign rom[13'h0a9c] = 1;
    assign rom[13'h0a9d] = 1;
    assign rom[13'h0a9e] = 1;
    assign rom[13'h0a9f] = 0;
    assign rom[13'h0aa0] = 0;
    assign rom[13'h0aa1] = 0;
    assign rom[13'h0aa2] = 1;
    assign rom[13'h0aa3] = 1;
    assign rom[13'h0aa4] = 1;
    assign rom[13'h0aa5] = 0;
    assign rom[13'h0aa6] = 0;
    assign rom[13'h0aa7] = 0;
    assign rom[13'h0aa8] = 0;
    assign rom[13'h0aa9] = 1;
    assign rom[13'h0aaa] = 1;
    assign rom[13'h0aab] = 0;
    assign rom[13'h0aac] = 1;
    assign rom[13'h0aad] = 1;
    assign rom[13'h0aae] = 0;
    assign rom[13'h0aaf] = 0;
    assign rom[13'h0ab0] = 0;
    assign rom[13'h0ab1] = 0;
    assign rom[13'h0ab2] = 0;
    assign rom[13'h0ab3] = 0;
    assign rom[13'h0ab4] = 0;
    assign rom[13'h0ab5] = 0;
    assign rom[13'h0ab6] = 0;
    assign rom[13'h0ab7] = 0;
    assign rom[13'h0ab8] = 0;
    assign rom[13'h0ab9] = 0;
    assign rom[13'h0aba] = 0;
    assign rom[13'h0abb] = 0;
    assign rom[13'h0abc] = 0;
    assign rom[13'h0abd] = 0;
    assign rom[13'h0abe] = 0;
    assign rom[13'h0abf] = 0;
    assign rom[13'h0ac0] = 0;
    assign rom[13'h0ac1] = 0;
    assign rom[13'h0ac2] = 0;
    assign rom[13'h0ac3] = 0;
    assign rom[13'h0ac4] = 0;
    assign rom[13'h0ac5] = 0;
    assign rom[13'h0ac6] = 0;
    assign rom[13'h0ac7] = 0;
    assign rom[13'h0ac8] = 0;
    assign rom[13'h0ac9] = 0;
    assign rom[13'h0aca] = 0;
    assign rom[13'h0acb] = 1;
    assign rom[13'h0acc] = 1;
    assign rom[13'h0acd] = 0;
    assign rom[13'h0ace] = 0;
    assign rom[13'h0acf] = 0;
    assign rom[13'h0ad0] = 0;
    assign rom[13'h0ad1] = 0;
    assign rom[13'h0ad2] = 0;
    assign rom[13'h0ad3] = 1;
    assign rom[13'h0ad4] = 1;
    assign rom[13'h0ad5] = 0;
    assign rom[13'h0ad6] = 0;
    assign rom[13'h0ad7] = 0;
    assign rom[13'h0ad8] = 0;
    assign rom[13'h0ad9] = 1;
    assign rom[13'h0ada] = 1;
    assign rom[13'h0adb] = 1;
    assign rom[13'h0adc] = 1;
    assign rom[13'h0add] = 1;
    assign rom[13'h0ade] = 1;
    assign rom[13'h0adf] = 0;
    assign rom[13'h0ae0] = 0;
    assign rom[13'h0ae1] = 0;
    assign rom[13'h0ae2] = 0;
    assign rom[13'h0ae3] = 1;
    assign rom[13'h0ae4] = 1;
    assign rom[13'h0ae5] = 0;
    assign rom[13'h0ae6] = 0;
    assign rom[13'h0ae7] = 0;
    assign rom[13'h0ae8] = 0;
    assign rom[13'h0ae9] = 0;
    assign rom[13'h0aea] = 0;
    assign rom[13'h0aeb] = 1;
    assign rom[13'h0aec] = 1;
    assign rom[13'h0aed] = 0;
    assign rom[13'h0aee] = 0;
    assign rom[13'h0aef] = 0;
    assign rom[13'h0af0] = 0;
    assign rom[13'h0af1] = 0;
    assign rom[13'h0af2] = 0;
    assign rom[13'h0af3] = 0;
    assign rom[13'h0af4] = 0;
    assign rom[13'h0af5] = 0;
    assign rom[13'h0af6] = 0;
    assign rom[13'h0af7] = 0;
    assign rom[13'h0af8] = 0;
    assign rom[13'h0af9] = 0;
    assign rom[13'h0afa] = 0;
    assign rom[13'h0afb] = 0;
    assign rom[13'h0afc] = 0;
    assign rom[13'h0afd] = 0;
    assign rom[13'h0afe] = 0;
    assign rom[13'h0aff] = 0;
    assign rom[13'h0b00] = 0;
    assign rom[13'h0b01] = 0;
    assign rom[13'h0b02] = 0;
    assign rom[13'h0b03] = 0;
    assign rom[13'h0b04] = 0;
    assign rom[13'h0b05] = 0;
    assign rom[13'h0b06] = 0;
    assign rom[13'h0b07] = 0;
    assign rom[13'h0b08] = 0;
    assign rom[13'h0b09] = 0;
    assign rom[13'h0b0a] = 0;
    assign rom[13'h0b0b] = 0;
    assign rom[13'h0b0c] = 0;
    assign rom[13'h0b0d] = 0;
    assign rom[13'h0b0e] = 0;
    assign rom[13'h0b0f] = 0;
    assign rom[13'h0b10] = 0;
    assign rom[13'h0b11] = 0;
    assign rom[13'h0b12] = 0;
    assign rom[13'h0b13] = 0;
    assign rom[13'h0b14] = 0;
    assign rom[13'h0b15] = 0;
    assign rom[13'h0b16] = 0;
    assign rom[13'h0b17] = 0;
    assign rom[13'h0b18] = 0;
    assign rom[13'h0b19] = 0;
    assign rom[13'h0b1a] = 0;
    assign rom[13'h0b1b] = 0;
    assign rom[13'h0b1c] = 0;
    assign rom[13'h0b1d] = 0;
    assign rom[13'h0b1e] = 0;
    assign rom[13'h0b1f] = 0;
    assign rom[13'h0b20] = 0;
    assign rom[13'h0b21] = 0;
    assign rom[13'h0b22] = 0;
    assign rom[13'h0b23] = 0;
    assign rom[13'h0b24] = 0;
    assign rom[13'h0b25] = 0;
    assign rom[13'h0b26] = 0;
    assign rom[13'h0b27] = 0;
    assign rom[13'h0b28] = 0;
    assign rom[13'h0b29] = 0;
    assign rom[13'h0b2a] = 0;
    assign rom[13'h0b2b] = 1;
    assign rom[13'h0b2c] = 1;
    assign rom[13'h0b2d] = 0;
    assign rom[13'h0b2e] = 0;
    assign rom[13'h0b2f] = 0;
    assign rom[13'h0b30] = 0;
    assign rom[13'h0b31] = 0;
    assign rom[13'h0b32] = 0;
    assign rom[13'h0b33] = 1;
    assign rom[13'h0b34] = 1;
    assign rom[13'h0b35] = 0;
    assign rom[13'h0b36] = 0;
    assign rom[13'h0b37] = 0;
    assign rom[13'h0b38] = 0;
    assign rom[13'h0b39] = 0;
    assign rom[13'h0b3a] = 0;
    assign rom[13'h0b3b] = 1;
    assign rom[13'h0b3c] = 0;
    assign rom[13'h0b3d] = 0;
    assign rom[13'h0b3e] = 0;
    assign rom[13'h0b3f] = 0;
    assign rom[13'h0b40] = 0;
    assign rom[13'h0b41] = 0;
    assign rom[13'h0b42] = 0;
    assign rom[13'h0b43] = 0;
    assign rom[13'h0b44] = 0;
    assign rom[13'h0b45] = 0;
    assign rom[13'h0b46] = 0;
    assign rom[13'h0b47] = 0;
    assign rom[13'h0b48] = 0;
    assign rom[13'h0b49] = 0;
    assign rom[13'h0b4a] = 0;
    assign rom[13'h0b4b] = 0;
    assign rom[13'h0b4c] = 0;
    assign rom[13'h0b4d] = 0;
    assign rom[13'h0b4e] = 0;
    assign rom[13'h0b4f] = 0;
    assign rom[13'h0b50] = 0;
    assign rom[13'h0b51] = 0;
    assign rom[13'h0b52] = 0;
    assign rom[13'h0b53] = 0;
    assign rom[13'h0b54] = 0;
    assign rom[13'h0b55] = 0;
    assign rom[13'h0b56] = 0;
    assign rom[13'h0b57] = 0;
    assign rom[13'h0b58] = 0;
    assign rom[13'h0b59] = 1;
    assign rom[13'h0b5a] = 1;
    assign rom[13'h0b5b] = 1;
    assign rom[13'h0b5c] = 1;
    assign rom[13'h0b5d] = 1;
    assign rom[13'h0b5e] = 1;
    assign rom[13'h0b5f] = 0;
    assign rom[13'h0b60] = 0;
    assign rom[13'h0b61] = 0;
    assign rom[13'h0b62] = 0;
    assign rom[13'h0b63] = 0;
    assign rom[13'h0b64] = 0;
    assign rom[13'h0b65] = 0;
    assign rom[13'h0b66] = 0;
    assign rom[13'h0b67] = 0;
    assign rom[13'h0b68] = 0;
    assign rom[13'h0b69] = 0;
    assign rom[13'h0b6a] = 0;
    assign rom[13'h0b6b] = 0;
    assign rom[13'h0b6c] = 0;
    assign rom[13'h0b6d] = 0;
    assign rom[13'h0b6e] = 0;
    assign rom[13'h0b6f] = 0;
    assign rom[13'h0b70] = 0;
    assign rom[13'h0b71] = 0;
    assign rom[13'h0b72] = 0;
    assign rom[13'h0b73] = 0;
    assign rom[13'h0b74] = 0;
    assign rom[13'h0b75] = 0;
    assign rom[13'h0b76] = 0;
    assign rom[13'h0b77] = 0;
    assign rom[13'h0b78] = 0;
    assign rom[13'h0b79] = 0;
    assign rom[13'h0b7a] = 0;
    assign rom[13'h0b7b] = 0;
    assign rom[13'h0b7c] = 0;
    assign rom[13'h0b7d] = 0;
    assign rom[13'h0b7e] = 0;
    assign rom[13'h0b7f] = 0;
    assign rom[13'h0b80] = 0;
    assign rom[13'h0b81] = 0;
    assign rom[13'h0b82] = 0;
    assign rom[13'h0b83] = 0;
    assign rom[13'h0b84] = 0;
    assign rom[13'h0b85] = 0;
    assign rom[13'h0b86] = 0;
    assign rom[13'h0b87] = 0;
    assign rom[13'h0b88] = 0;
    assign rom[13'h0b89] = 0;
    assign rom[13'h0b8a] = 0;
    assign rom[13'h0b8b] = 0;
    assign rom[13'h0b8c] = 0;
    assign rom[13'h0b8d] = 0;
    assign rom[13'h0b8e] = 0;
    assign rom[13'h0b8f] = 0;
    assign rom[13'h0b90] = 0;
    assign rom[13'h0b91] = 0;
    assign rom[13'h0b92] = 0;
    assign rom[13'h0b93] = 0;
    assign rom[13'h0b94] = 0;
    assign rom[13'h0b95] = 0;
    assign rom[13'h0b96] = 0;
    assign rom[13'h0b97] = 0;
    assign rom[13'h0b98] = 0;
    assign rom[13'h0b99] = 0;
    assign rom[13'h0b9a] = 0;
    assign rom[13'h0b9b] = 0;
    assign rom[13'h0b9c] = 0;
    assign rom[13'h0b9d] = 0;
    assign rom[13'h0b9e] = 0;
    assign rom[13'h0b9f] = 0;
    assign rom[13'h0ba0] = 0;
    assign rom[13'h0ba1] = 0;
    assign rom[13'h0ba2] = 0;
    assign rom[13'h0ba3] = 0;
    assign rom[13'h0ba4] = 0;
    assign rom[13'h0ba5] = 0;
    assign rom[13'h0ba6] = 0;
    assign rom[13'h0ba7] = 0;
    assign rom[13'h0ba8] = 0;
    assign rom[13'h0ba9] = 0;
    assign rom[13'h0baa] = 0;
    assign rom[13'h0bab] = 1;
    assign rom[13'h0bac] = 1;
    assign rom[13'h0bad] = 0;
    assign rom[13'h0bae] = 0;
    assign rom[13'h0baf] = 0;
    assign rom[13'h0bb0] = 0;
    assign rom[13'h0bb1] = 0;
    assign rom[13'h0bb2] = 0;
    assign rom[13'h0bb3] = 1;
    assign rom[13'h0bb4] = 1;
    assign rom[13'h0bb5] = 0;
    assign rom[13'h0bb6] = 0;
    assign rom[13'h0bb7] = 0;
    assign rom[13'h0bb8] = 0;
    assign rom[13'h0bb9] = 0;
    assign rom[13'h0bba] = 0;
    assign rom[13'h0bbb] = 0;
    assign rom[13'h0bbc] = 0;
    assign rom[13'h0bbd] = 0;
    assign rom[13'h0bbe] = 0;
    assign rom[13'h0bbf] = 0;
    assign rom[13'h0bc0] = 0;
    assign rom[13'h0bc1] = 0;
    assign rom[13'h0bc2] = 0;
    assign rom[13'h0bc3] = 0;
    assign rom[13'h0bc4] = 0;
    assign rom[13'h0bc5] = 0;
    assign rom[13'h0bc6] = 1;
    assign rom[13'h0bc7] = 0;
    assign rom[13'h0bc8] = 0;
    assign rom[13'h0bc9] = 0;
    assign rom[13'h0bca] = 0;
    assign rom[13'h0bcb] = 0;
    assign rom[13'h0bcc] = 0;
    assign rom[13'h0bcd] = 1;
    assign rom[13'h0bce] = 1;
    assign rom[13'h0bcf] = 0;
    assign rom[13'h0bd0] = 0;
    assign rom[13'h0bd1] = 0;
    assign rom[13'h0bd2] = 0;
    assign rom[13'h0bd3] = 0;
    assign rom[13'h0bd4] = 1;
    assign rom[13'h0bd5] = 1;
    assign rom[13'h0bd6] = 0;
    assign rom[13'h0bd7] = 0;
    assign rom[13'h0bd8] = 0;
    assign rom[13'h0bd9] = 0;
    assign rom[13'h0bda] = 0;
    assign rom[13'h0bdb] = 1;
    assign rom[13'h0bdc] = 1;
    assign rom[13'h0bdd] = 0;
    assign rom[13'h0bde] = 0;
    assign rom[13'h0bdf] = 0;
    assign rom[13'h0be0] = 0;
    assign rom[13'h0be1] = 0;
    assign rom[13'h0be2] = 1;
    assign rom[13'h0be3] = 1;
    assign rom[13'h0be4] = 0;
    assign rom[13'h0be5] = 0;
    assign rom[13'h0be6] = 0;
    assign rom[13'h0be7] = 0;
    assign rom[13'h0be8] = 0;
    assign rom[13'h0be9] = 1;
    assign rom[13'h0bea] = 1;
    assign rom[13'h0beb] = 0;
    assign rom[13'h0bec] = 0;
    assign rom[13'h0bed] = 0;
    assign rom[13'h0bee] = 0;
    assign rom[13'h0bef] = 0;
    assign rom[13'h0bf0] = 0;
    assign rom[13'h0bf1] = 1;
    assign rom[13'h0bf2] = 0;
    assign rom[13'h0bf3] = 0;
    assign rom[13'h0bf4] = 0;
    assign rom[13'h0bf5] = 0;
    assign rom[13'h0bf6] = 0;
    assign rom[13'h0bf7] = 0;
    assign rom[13'h0bf8] = 0;
    assign rom[13'h0bf9] = 0;
    assign rom[13'h0bfa] = 0;
    assign rom[13'h0bfb] = 0;
    assign rom[13'h0bfc] = 0;
    assign rom[13'h0bfd] = 0;
    assign rom[13'h0bfe] = 0;
    assign rom[13'h0bff] = 0;
    assign rom[13'h0c00] = 0;
    assign rom[13'h0c01] = 0;
    assign rom[13'h0c02] = 1;
    assign rom[13'h0c03] = 1;
    assign rom[13'h0c04] = 1;
    assign rom[13'h0c05] = 1;
    assign rom[13'h0c06] = 0;
    assign rom[13'h0c07] = 0;
    assign rom[13'h0c08] = 0;
    assign rom[13'h0c09] = 1;
    assign rom[13'h0c0a] = 1;
    assign rom[13'h0c0b] = 0;
    assign rom[13'h0c0c] = 0;
    assign rom[13'h0c0d] = 1;
    assign rom[13'h0c0e] = 1;
    assign rom[13'h0c0f] = 0;
    assign rom[13'h0c10] = 0;
    assign rom[13'h0c11] = 1;
    assign rom[13'h0c12] = 1;
    assign rom[13'h0c13] = 0;
    assign rom[13'h0c14] = 1;
    assign rom[13'h0c15] = 1;
    assign rom[13'h0c16] = 1;
    assign rom[13'h0c17] = 0;
    assign rom[13'h0c18] = 0;
    assign rom[13'h0c19] = 1;
    assign rom[13'h0c1a] = 1;
    assign rom[13'h0c1b] = 1;
    assign rom[13'h0c1c] = 0;
    assign rom[13'h0c1d] = 1;
    assign rom[13'h0c1e] = 1;
    assign rom[13'h0c1f] = 0;
    assign rom[13'h0c20] = 0;
    assign rom[13'h0c21] = 1;
    assign rom[13'h0c22] = 1;
    assign rom[13'h0c23] = 0;
    assign rom[13'h0c24] = 0;
    assign rom[13'h0c25] = 1;
    assign rom[13'h0c26] = 1;
    assign rom[13'h0c27] = 0;
    assign rom[13'h0c28] = 0;
    assign rom[13'h0c29] = 1;
    assign rom[13'h0c2a] = 1;
    assign rom[13'h0c2b] = 0;
    assign rom[13'h0c2c] = 0;
    assign rom[13'h0c2d] = 1;
    assign rom[13'h0c2e] = 1;
    assign rom[13'h0c2f] = 0;
    assign rom[13'h0c30] = 0;
    assign rom[13'h0c31] = 0;
    assign rom[13'h0c32] = 1;
    assign rom[13'h0c33] = 1;
    assign rom[13'h0c34] = 1;
    assign rom[13'h0c35] = 1;
    assign rom[13'h0c36] = 0;
    assign rom[13'h0c37] = 0;
    assign rom[13'h0c38] = 0;
    assign rom[13'h0c39] = 0;
    assign rom[13'h0c3a] = 0;
    assign rom[13'h0c3b] = 0;
    assign rom[13'h0c3c] = 0;
    assign rom[13'h0c3d] = 0;
    assign rom[13'h0c3e] = 0;
    assign rom[13'h0c3f] = 0;
    assign rom[13'h0c40] = 0;
    assign rom[13'h0c41] = 0;
    assign rom[13'h0c42] = 0;
    assign rom[13'h0c43] = 1;
    assign rom[13'h0c44] = 1;
    assign rom[13'h0c45] = 0;
    assign rom[13'h0c46] = 0;
    assign rom[13'h0c47] = 0;
    assign rom[13'h0c48] = 0;
    assign rom[13'h0c49] = 0;
    assign rom[13'h0c4a] = 0;
    assign rom[13'h0c4b] = 1;
    assign rom[13'h0c4c] = 1;
    assign rom[13'h0c4d] = 0;
    assign rom[13'h0c4e] = 0;
    assign rom[13'h0c4f] = 0;
    assign rom[13'h0c50] = 0;
    assign rom[13'h0c51] = 0;
    assign rom[13'h0c52] = 1;
    assign rom[13'h0c53] = 1;
    assign rom[13'h0c54] = 1;
    assign rom[13'h0c55] = 0;
    assign rom[13'h0c56] = 0;
    assign rom[13'h0c57] = 0;
    assign rom[13'h0c58] = 0;
    assign rom[13'h0c59] = 0;
    assign rom[13'h0c5a] = 0;
    assign rom[13'h0c5b] = 1;
    assign rom[13'h0c5c] = 1;
    assign rom[13'h0c5d] = 0;
    assign rom[13'h0c5e] = 0;
    assign rom[13'h0c5f] = 0;
    assign rom[13'h0c60] = 0;
    assign rom[13'h0c61] = 0;
    assign rom[13'h0c62] = 0;
    assign rom[13'h0c63] = 1;
    assign rom[13'h0c64] = 1;
    assign rom[13'h0c65] = 0;
    assign rom[13'h0c66] = 0;
    assign rom[13'h0c67] = 0;
    assign rom[13'h0c68] = 0;
    assign rom[13'h0c69] = 0;
    assign rom[13'h0c6a] = 0;
    assign rom[13'h0c6b] = 1;
    assign rom[13'h0c6c] = 1;
    assign rom[13'h0c6d] = 0;
    assign rom[13'h0c6e] = 0;
    assign rom[13'h0c6f] = 0;
    assign rom[13'h0c70] = 0;
    assign rom[13'h0c71] = 0;
    assign rom[13'h0c72] = 1;
    assign rom[13'h0c73] = 1;
    assign rom[13'h0c74] = 1;
    assign rom[13'h0c75] = 1;
    assign rom[13'h0c76] = 0;
    assign rom[13'h0c77] = 0;
    assign rom[13'h0c78] = 0;
    assign rom[13'h0c79] = 0;
    assign rom[13'h0c7a] = 0;
    assign rom[13'h0c7b] = 0;
    assign rom[13'h0c7c] = 0;
    assign rom[13'h0c7d] = 0;
    assign rom[13'h0c7e] = 0;
    assign rom[13'h0c7f] = 0;
    assign rom[13'h0c80] = 0;
    assign rom[13'h0c81] = 1;
    assign rom[13'h0c82] = 1;
    assign rom[13'h0c83] = 1;
    assign rom[13'h0c84] = 1;
    assign rom[13'h0c85] = 1;
    assign rom[13'h0c86] = 0;
    assign rom[13'h0c87] = 0;
    assign rom[13'h0c88] = 0;
    assign rom[13'h0c89] = 0;
    assign rom[13'h0c8a] = 0;
    assign rom[13'h0c8b] = 0;
    assign rom[13'h0c8c] = 0;
    assign rom[13'h0c8d] = 1;
    assign rom[13'h0c8e] = 1;
    assign rom[13'h0c8f] = 0;
    assign rom[13'h0c90] = 0;
    assign rom[13'h0c91] = 0;
    assign rom[13'h0c92] = 0;
    assign rom[13'h0c93] = 0;
    assign rom[13'h0c94] = 0;
    assign rom[13'h0c95] = 1;
    assign rom[13'h0c96] = 1;
    assign rom[13'h0c97] = 0;
    assign rom[13'h0c98] = 0;
    assign rom[13'h0c99] = 0;
    assign rom[13'h0c9a] = 1;
    assign rom[13'h0c9b] = 1;
    assign rom[13'h0c9c] = 1;
    assign rom[13'h0c9d] = 1;
    assign rom[13'h0c9e] = 0;
    assign rom[13'h0c9f] = 0;
    assign rom[13'h0ca0] = 0;
    assign rom[13'h0ca1] = 1;
    assign rom[13'h0ca2] = 1;
    assign rom[13'h0ca3] = 0;
    assign rom[13'h0ca4] = 0;
    assign rom[13'h0ca5] = 0;
    assign rom[13'h0ca6] = 0;
    assign rom[13'h0ca7] = 0;
    assign rom[13'h0ca8] = 0;
    assign rom[13'h0ca9] = 1;
    assign rom[13'h0caa] = 1;
    assign rom[13'h0cab] = 0;
    assign rom[13'h0cac] = 0;
    assign rom[13'h0cad] = 0;
    assign rom[13'h0cae] = 0;
    assign rom[13'h0caf] = 0;
    assign rom[13'h0cb0] = 0;
    assign rom[13'h0cb1] = 1;
    assign rom[13'h0cb2] = 1;
    assign rom[13'h0cb3] = 1;
    assign rom[13'h0cb4] = 1;
    assign rom[13'h0cb5] = 1;
    assign rom[13'h0cb6] = 0;
    assign rom[13'h0cb7] = 0;
    assign rom[13'h0cb8] = 0;
    assign rom[13'h0cb9] = 0;
    assign rom[13'h0cba] = 0;
    assign rom[13'h0cbb] = 0;
    assign rom[13'h0cbc] = 0;
    assign rom[13'h0cbd] = 0;
    assign rom[13'h0cbe] = 0;
    assign rom[13'h0cbf] = 0;
    assign rom[13'h0cc0] = 0;
    assign rom[13'h0cc1] = 1;
    assign rom[13'h0cc2] = 1;
    assign rom[13'h0cc3] = 1;
    assign rom[13'h0cc4] = 1;
    assign rom[13'h0cc5] = 1;
    assign rom[13'h0cc6] = 0;
    assign rom[13'h0cc7] = 0;
    assign rom[13'h0cc8] = 0;
    assign rom[13'h0cc9] = 0;
    assign rom[13'h0cca] = 0;
    assign rom[13'h0ccb] = 0;
    assign rom[13'h0ccc] = 0;
    assign rom[13'h0ccd] = 1;
    assign rom[13'h0cce] = 1;
    assign rom[13'h0ccf] = 0;
    assign rom[13'h0cd0] = 0;
    assign rom[13'h0cd1] = 0;
    assign rom[13'h0cd2] = 0;
    assign rom[13'h0cd3] = 0;
    assign rom[13'h0cd4] = 0;
    assign rom[13'h0cd5] = 1;
    assign rom[13'h0cd6] = 1;
    assign rom[13'h0cd7] = 0;
    assign rom[13'h0cd8] = 0;
    assign rom[13'h0cd9] = 0;
    assign rom[13'h0cda] = 1;
    assign rom[13'h0cdb] = 1;
    assign rom[13'h0cdc] = 1;
    assign rom[13'h0cdd] = 1;
    assign rom[13'h0cde] = 0;
    assign rom[13'h0cdf] = 0;
    assign rom[13'h0ce0] = 0;
    assign rom[13'h0ce1] = 0;
    assign rom[13'h0ce2] = 0;
    assign rom[13'h0ce3] = 0;
    assign rom[13'h0ce4] = 0;
    assign rom[13'h0ce5] = 1;
    assign rom[13'h0ce6] = 1;
    assign rom[13'h0ce7] = 0;
    assign rom[13'h0ce8] = 0;
    assign rom[13'h0ce9] = 0;
    assign rom[13'h0cea] = 0;
    assign rom[13'h0ceb] = 0;
    assign rom[13'h0cec] = 0;
    assign rom[13'h0ced] = 1;
    assign rom[13'h0cee] = 1;
    assign rom[13'h0cef] = 0;
    assign rom[13'h0cf0] = 0;
    assign rom[13'h0cf1] = 1;
    assign rom[13'h0cf2] = 1;
    assign rom[13'h0cf3] = 1;
    assign rom[13'h0cf4] = 1;
    assign rom[13'h0cf5] = 1;
    assign rom[13'h0cf6] = 0;
    assign rom[13'h0cf7] = 0;
    assign rom[13'h0cf8] = 0;
    assign rom[13'h0cf9] = 0;
    assign rom[13'h0cfa] = 0;
    assign rom[13'h0cfb] = 0;
    assign rom[13'h0cfc] = 0;
    assign rom[13'h0cfd] = 0;
    assign rom[13'h0cfe] = 0;
    assign rom[13'h0cff] = 0;
    assign rom[13'h0d00] = 0;
    assign rom[13'h0d01] = 1;
    assign rom[13'h0d02] = 1;
    assign rom[13'h0d03] = 0;
    assign rom[13'h0d04] = 0;
    assign rom[13'h0d05] = 1;
    assign rom[13'h0d06] = 1;
    assign rom[13'h0d07] = 0;
    assign rom[13'h0d08] = 0;
    assign rom[13'h0d09] = 1;
    assign rom[13'h0d0a] = 1;
    assign rom[13'h0d0b] = 0;
    assign rom[13'h0d0c] = 0;
    assign rom[13'h0d0d] = 1;
    assign rom[13'h0d0e] = 1;
    assign rom[13'h0d0f] = 0;
    assign rom[13'h0d10] = 0;
    assign rom[13'h0d11] = 1;
    assign rom[13'h0d12] = 1;
    assign rom[13'h0d13] = 0;
    assign rom[13'h0d14] = 0;
    assign rom[13'h0d15] = 1;
    assign rom[13'h0d16] = 1;
    assign rom[13'h0d17] = 0;
    assign rom[13'h0d18] = 0;
    assign rom[13'h0d19] = 1;
    assign rom[13'h0d1a] = 1;
    assign rom[13'h0d1b] = 1;
    assign rom[13'h0d1c] = 1;
    assign rom[13'h0d1d] = 1;
    assign rom[13'h0d1e] = 1;
    assign rom[13'h0d1f] = 0;
    assign rom[13'h0d20] = 0;
    assign rom[13'h0d21] = 0;
    assign rom[13'h0d22] = 0;
    assign rom[13'h0d23] = 0;
    assign rom[13'h0d24] = 0;
    assign rom[13'h0d25] = 1;
    assign rom[13'h0d26] = 1;
    assign rom[13'h0d27] = 0;
    assign rom[13'h0d28] = 0;
    assign rom[13'h0d29] = 0;
    assign rom[13'h0d2a] = 0;
    assign rom[13'h0d2b] = 0;
    assign rom[13'h0d2c] = 0;
    assign rom[13'h0d2d] = 1;
    assign rom[13'h0d2e] = 1;
    assign rom[13'h0d2f] = 0;
    assign rom[13'h0d30] = 0;
    assign rom[13'h0d31] = 0;
    assign rom[13'h0d32] = 0;
    assign rom[13'h0d33] = 0;
    assign rom[13'h0d34] = 0;
    assign rom[13'h0d35] = 1;
    assign rom[13'h0d36] = 1;
    assign rom[13'h0d37] = 0;
    assign rom[13'h0d38] = 0;
    assign rom[13'h0d39] = 0;
    assign rom[13'h0d3a] = 0;
    assign rom[13'h0d3b] = 0;
    assign rom[13'h0d3c] = 0;
    assign rom[13'h0d3d] = 0;
    assign rom[13'h0d3e] = 0;
    assign rom[13'h0d3f] = 0;
    assign rom[13'h0d40] = 0;
    assign rom[13'h0d41] = 1;
    assign rom[13'h0d42] = 1;
    assign rom[13'h0d43] = 1;
    assign rom[13'h0d44] = 1;
    assign rom[13'h0d45] = 1;
    assign rom[13'h0d46] = 1;
    assign rom[13'h0d47] = 0;
    assign rom[13'h0d48] = 0;
    assign rom[13'h0d49] = 1;
    assign rom[13'h0d4a] = 1;
    assign rom[13'h0d4b] = 0;
    assign rom[13'h0d4c] = 0;
    assign rom[13'h0d4d] = 0;
    assign rom[13'h0d4e] = 0;
    assign rom[13'h0d4f] = 0;
    assign rom[13'h0d50] = 0;
    assign rom[13'h0d51] = 1;
    assign rom[13'h0d52] = 1;
    assign rom[13'h0d53] = 0;
    assign rom[13'h0d54] = 0;
    assign rom[13'h0d55] = 0;
    assign rom[13'h0d56] = 0;
    assign rom[13'h0d57] = 0;
    assign rom[13'h0d58] = 0;
    assign rom[13'h0d59] = 1;
    assign rom[13'h0d5a] = 1;
    assign rom[13'h0d5b] = 1;
    assign rom[13'h0d5c] = 1;
    assign rom[13'h0d5d] = 1;
    assign rom[13'h0d5e] = 0;
    assign rom[13'h0d5f] = 0;
    assign rom[13'h0d60] = 0;
    assign rom[13'h0d61] = 0;
    assign rom[13'h0d62] = 0;
    assign rom[13'h0d63] = 0;
    assign rom[13'h0d64] = 0;
    assign rom[13'h0d65] = 1;
    assign rom[13'h0d66] = 1;
    assign rom[13'h0d67] = 0;
    assign rom[13'h0d68] = 0;
    assign rom[13'h0d69] = 0;
    assign rom[13'h0d6a] = 0;
    assign rom[13'h0d6b] = 0;
    assign rom[13'h0d6c] = 0;
    assign rom[13'h0d6d] = 1;
    assign rom[13'h0d6e] = 1;
    assign rom[13'h0d6f] = 0;
    assign rom[13'h0d70] = 0;
    assign rom[13'h0d71] = 1;
    assign rom[13'h0d72] = 1;
    assign rom[13'h0d73] = 1;
    assign rom[13'h0d74] = 1;
    assign rom[13'h0d75] = 1;
    assign rom[13'h0d76] = 0;
    assign rom[13'h0d77] = 0;
    assign rom[13'h0d78] = 0;
    assign rom[13'h0d79] = 0;
    assign rom[13'h0d7a] = 0;
    assign rom[13'h0d7b] = 0;
    assign rom[13'h0d7c] = 0;
    assign rom[13'h0d7d] = 0;
    assign rom[13'h0d7e] = 0;
    assign rom[13'h0d7f] = 0;
    assign rom[13'h0d80] = 0;
    assign rom[13'h0d81] = 0;
    assign rom[13'h0d82] = 1;
    assign rom[13'h0d83] = 1;
    assign rom[13'h0d84] = 1;
    assign rom[13'h0d85] = 1;
    assign rom[13'h0d86] = 0;
    assign rom[13'h0d87] = 0;
    assign rom[13'h0d88] = 0;
    assign rom[13'h0d89] = 1;
    assign rom[13'h0d8a] = 1;
    assign rom[13'h0d8b] = 0;
    assign rom[13'h0d8c] = 0;
    assign rom[13'h0d8d] = 0;
    assign rom[13'h0d8e] = 0;
    assign rom[13'h0d8f] = 0;
    assign rom[13'h0d90] = 0;
    assign rom[13'h0d91] = 1;
    assign rom[13'h0d92] = 1;
    assign rom[13'h0d93] = 0;
    assign rom[13'h0d94] = 0;
    assign rom[13'h0d95] = 0;
    assign rom[13'h0d96] = 0;
    assign rom[13'h0d97] = 0;
    assign rom[13'h0d98] = 0;
    assign rom[13'h0d99] = 1;
    assign rom[13'h0d9a] = 1;
    assign rom[13'h0d9b] = 1;
    assign rom[13'h0d9c] = 1;
    assign rom[13'h0d9d] = 1;
    assign rom[13'h0d9e] = 0;
    assign rom[13'h0d9f] = 0;
    assign rom[13'h0da0] = 0;
    assign rom[13'h0da1] = 1;
    assign rom[13'h0da2] = 1;
    assign rom[13'h0da3] = 0;
    assign rom[13'h0da4] = 0;
    assign rom[13'h0da5] = 1;
    assign rom[13'h0da6] = 1;
    assign rom[13'h0da7] = 0;
    assign rom[13'h0da8] = 0;
    assign rom[13'h0da9] = 1;
    assign rom[13'h0daa] = 1;
    assign rom[13'h0dab] = 0;
    assign rom[13'h0dac] = 0;
    assign rom[13'h0dad] = 1;
    assign rom[13'h0dae] = 1;
    assign rom[13'h0daf] = 0;
    assign rom[13'h0db0] = 0;
    assign rom[13'h0db1] = 0;
    assign rom[13'h0db2] = 1;
    assign rom[13'h0db3] = 1;
    assign rom[13'h0db4] = 1;
    assign rom[13'h0db5] = 1;
    assign rom[13'h0db6] = 0;
    assign rom[13'h0db7] = 0;
    assign rom[13'h0db8] = 0;
    assign rom[13'h0db9] = 0;
    assign rom[13'h0dba] = 0;
    assign rom[13'h0dbb] = 0;
    assign rom[13'h0dbc] = 0;
    assign rom[13'h0dbd] = 0;
    assign rom[13'h0dbe] = 0;
    assign rom[13'h0dbf] = 0;
    assign rom[13'h0dc0] = 0;
    assign rom[13'h0dc1] = 1;
    assign rom[13'h0dc2] = 1;
    assign rom[13'h0dc3] = 1;
    assign rom[13'h0dc4] = 1;
    assign rom[13'h0dc5] = 1;
    assign rom[13'h0dc6] = 1;
    assign rom[13'h0dc7] = 0;
    assign rom[13'h0dc8] = 0;
    assign rom[13'h0dc9] = 0;
    assign rom[13'h0dca] = 0;
    assign rom[13'h0dcb] = 0;
    assign rom[13'h0dcc] = 0;
    assign rom[13'h0dcd] = 1;
    assign rom[13'h0dce] = 1;
    assign rom[13'h0dcf] = 0;
    assign rom[13'h0dd0] = 0;
    assign rom[13'h0dd1] = 0;
    assign rom[13'h0dd2] = 0;
    assign rom[13'h0dd3] = 0;
    assign rom[13'h0dd4] = 1;
    assign rom[13'h0dd5] = 1;
    assign rom[13'h0dd6] = 0;
    assign rom[13'h0dd7] = 0;
    assign rom[13'h0dd8] = 0;
    assign rom[13'h0dd9] = 0;
    assign rom[13'h0dda] = 0;
    assign rom[13'h0ddb] = 1;
    assign rom[13'h0ddc] = 1;
    assign rom[13'h0ddd] = 0;
    assign rom[13'h0dde] = 0;
    assign rom[13'h0ddf] = 0;
    assign rom[13'h0de0] = 0;
    assign rom[13'h0de1] = 0;
    assign rom[13'h0de2] = 0;
    assign rom[13'h0de3] = 1;
    assign rom[13'h0de4] = 1;
    assign rom[13'h0de5] = 0;
    assign rom[13'h0de6] = 0;
    assign rom[13'h0de7] = 0;
    assign rom[13'h0de8] = 0;
    assign rom[13'h0de9] = 0;
    assign rom[13'h0dea] = 0;
    assign rom[13'h0deb] = 1;
    assign rom[13'h0dec] = 1;
    assign rom[13'h0ded] = 0;
    assign rom[13'h0dee] = 0;
    assign rom[13'h0def] = 0;
    assign rom[13'h0df0] = 0;
    assign rom[13'h0df1] = 0;
    assign rom[13'h0df2] = 0;
    assign rom[13'h0df3] = 1;
    assign rom[13'h0df4] = 1;
    assign rom[13'h0df5] = 0;
    assign rom[13'h0df6] = 0;
    assign rom[13'h0df7] = 0;
    assign rom[13'h0df8] = 0;
    assign rom[13'h0df9] = 0;
    assign rom[13'h0dfa] = 0;
    assign rom[13'h0dfb] = 0;
    assign rom[13'h0dfc] = 0;
    assign rom[13'h0dfd] = 0;
    assign rom[13'h0dfe] = 0;
    assign rom[13'h0dff] = 0;
    assign rom[13'h0e00] = 0;
    assign rom[13'h0e01] = 0;
    assign rom[13'h0e02] = 1;
    assign rom[13'h0e03] = 1;
    assign rom[13'h0e04] = 1;
    assign rom[13'h0e05] = 1;
    assign rom[13'h0e06] = 0;
    assign rom[13'h0e07] = 0;
    assign rom[13'h0e08] = 0;
    assign rom[13'h0e09] = 1;
    assign rom[13'h0e0a] = 1;
    assign rom[13'h0e0b] = 0;
    assign rom[13'h0e0c] = 0;
    assign rom[13'h0e0d] = 1;
    assign rom[13'h0e0e] = 1;
    assign rom[13'h0e0f] = 0;
    assign rom[13'h0e10] = 0;
    assign rom[13'h0e11] = 1;
    assign rom[13'h0e12] = 1;
    assign rom[13'h0e13] = 0;
    assign rom[13'h0e14] = 0;
    assign rom[13'h0e15] = 1;
    assign rom[13'h0e16] = 1;
    assign rom[13'h0e17] = 0;
    assign rom[13'h0e18] = 0;
    assign rom[13'h0e19] = 0;
    assign rom[13'h0e1a] = 1;
    assign rom[13'h0e1b] = 1;
    assign rom[13'h0e1c] = 1;
    assign rom[13'h0e1d] = 1;
    assign rom[13'h0e1e] = 0;
    assign rom[13'h0e1f] = 0;
    assign rom[13'h0e20] = 0;
    assign rom[13'h0e21] = 1;
    assign rom[13'h0e22] = 1;
    assign rom[13'h0e23] = 0;
    assign rom[13'h0e24] = 0;
    assign rom[13'h0e25] = 1;
    assign rom[13'h0e26] = 1;
    assign rom[13'h0e27] = 0;
    assign rom[13'h0e28] = 0;
    assign rom[13'h0e29] = 1;
    assign rom[13'h0e2a] = 1;
    assign rom[13'h0e2b] = 0;
    assign rom[13'h0e2c] = 0;
    assign rom[13'h0e2d] = 1;
    assign rom[13'h0e2e] = 1;
    assign rom[13'h0e2f] = 0;
    assign rom[13'h0e30] = 0;
    assign rom[13'h0e31] = 0;
    assign rom[13'h0e32] = 1;
    assign rom[13'h0e33] = 1;
    assign rom[13'h0e34] = 1;
    assign rom[13'h0e35] = 1;
    assign rom[13'h0e36] = 0;
    assign rom[13'h0e37] = 0;
    assign rom[13'h0e38] = 0;
    assign rom[13'h0e39] = 0;
    assign rom[13'h0e3a] = 0;
    assign rom[13'h0e3b] = 0;
    assign rom[13'h0e3c] = 0;
    assign rom[13'h0e3d] = 0;
    assign rom[13'h0e3e] = 0;
    assign rom[13'h0e3f] = 0;
    assign rom[13'h0e40] = 0;
    assign rom[13'h0e41] = 0;
    assign rom[13'h0e42] = 1;
    assign rom[13'h0e43] = 1;
    assign rom[13'h0e44] = 1;
    assign rom[13'h0e45] = 1;
    assign rom[13'h0e46] = 0;
    assign rom[13'h0e47] = 0;
    assign rom[13'h0e48] = 0;
    assign rom[13'h0e49] = 1;
    assign rom[13'h0e4a] = 1;
    assign rom[13'h0e4b] = 0;
    assign rom[13'h0e4c] = 0;
    assign rom[13'h0e4d] = 1;
    assign rom[13'h0e4e] = 1;
    assign rom[13'h0e4f] = 0;
    assign rom[13'h0e50] = 0;
    assign rom[13'h0e51] = 1;
    assign rom[13'h0e52] = 1;
    assign rom[13'h0e53] = 0;
    assign rom[13'h0e54] = 0;
    assign rom[13'h0e55] = 1;
    assign rom[13'h0e56] = 1;
    assign rom[13'h0e57] = 0;
    assign rom[13'h0e58] = 0;
    assign rom[13'h0e59] = 0;
    assign rom[13'h0e5a] = 1;
    assign rom[13'h0e5b] = 1;
    assign rom[13'h0e5c] = 1;
    assign rom[13'h0e5d] = 1;
    assign rom[13'h0e5e] = 1;
    assign rom[13'h0e5f] = 0;
    assign rom[13'h0e60] = 0;
    assign rom[13'h0e61] = 0;
    assign rom[13'h0e62] = 0;
    assign rom[13'h0e63] = 0;
    assign rom[13'h0e64] = 0;
    assign rom[13'h0e65] = 1;
    assign rom[13'h0e66] = 1;
    assign rom[13'h0e67] = 0;
    assign rom[13'h0e68] = 0;
    assign rom[13'h0e69] = 0;
    assign rom[13'h0e6a] = 0;
    assign rom[13'h0e6b] = 0;
    assign rom[13'h0e6c] = 0;
    assign rom[13'h0e6d] = 1;
    assign rom[13'h0e6e] = 1;
    assign rom[13'h0e6f] = 0;
    assign rom[13'h0e70] = 0;
    assign rom[13'h0e71] = 0;
    assign rom[13'h0e72] = 1;
    assign rom[13'h0e73] = 1;
    assign rom[13'h0e74] = 1;
    assign rom[13'h0e75] = 1;
    assign rom[13'h0e76] = 0;
    assign rom[13'h0e77] = 0;
    assign rom[13'h0e78] = 0;
    assign rom[13'h0e79] = 0;
    assign rom[13'h0e7a] = 0;
    assign rom[13'h0e7b] = 0;
    assign rom[13'h0e7c] = 0;
    assign rom[13'h0e7d] = 0;
    assign rom[13'h0e7e] = 0;
    assign rom[13'h0e7f] = 0;
    assign rom[13'h0e80] = 0;
    assign rom[13'h0e81] = 0;
    assign rom[13'h0e82] = 0;
    assign rom[13'h0e83] = 0;
    assign rom[13'h0e84] = 0;
    assign rom[13'h0e85] = 0;
    assign rom[13'h0e86] = 0;
    assign rom[13'h0e87] = 0;
    assign rom[13'h0e88] = 0;
    assign rom[13'h0e89] = 0;
    assign rom[13'h0e8a] = 0;
    assign rom[13'h0e8b] = 1;
    assign rom[13'h0e8c] = 1;
    assign rom[13'h0e8d] = 0;
    assign rom[13'h0e8e] = 0;
    assign rom[13'h0e8f] = 0;
    assign rom[13'h0e90] = 0;
    assign rom[13'h0e91] = 0;
    assign rom[13'h0e92] = 0;
    assign rom[13'h0e93] = 1;
    assign rom[13'h0e94] = 1;
    assign rom[13'h0e95] = 0;
    assign rom[13'h0e96] = 0;
    assign rom[13'h0e97] = 0;
    assign rom[13'h0e98] = 0;
    assign rom[13'h0e99] = 0;
    assign rom[13'h0e9a] = 0;
    assign rom[13'h0e9b] = 0;
    assign rom[13'h0e9c] = 0;
    assign rom[13'h0e9d] = 0;
    assign rom[13'h0e9e] = 0;
    assign rom[13'h0e9f] = 0;
    assign rom[13'h0ea0] = 0;
    assign rom[13'h0ea1] = 0;
    assign rom[13'h0ea2] = 0;
    assign rom[13'h0ea3] = 1;
    assign rom[13'h0ea4] = 1;
    assign rom[13'h0ea5] = 0;
    assign rom[13'h0ea6] = 0;
    assign rom[13'h0ea7] = 0;
    assign rom[13'h0ea8] = 0;
    assign rom[13'h0ea9] = 0;
    assign rom[13'h0eaa] = 0;
    assign rom[13'h0eab] = 1;
    assign rom[13'h0eac] = 1;
    assign rom[13'h0ead] = 0;
    assign rom[13'h0eae] = 0;
    assign rom[13'h0eaf] = 0;
    assign rom[13'h0eb0] = 0;
    assign rom[13'h0eb1] = 0;
    assign rom[13'h0eb2] = 0;
    assign rom[13'h0eb3] = 0;
    assign rom[13'h0eb4] = 0;
    assign rom[13'h0eb5] = 0;
    assign rom[13'h0eb6] = 0;
    assign rom[13'h0eb7] = 0;
    assign rom[13'h0eb8] = 0;
    assign rom[13'h0eb9] = 0;
    assign rom[13'h0eba] = 0;
    assign rom[13'h0ebb] = 0;
    assign rom[13'h0ebc] = 0;
    assign rom[13'h0ebd] = 0;
    assign rom[13'h0ebe] = 0;
    assign rom[13'h0ebf] = 0;
    assign rom[13'h0ec0] = 0;
    assign rom[13'h0ec1] = 0;
    assign rom[13'h0ec2] = 0;
    assign rom[13'h0ec3] = 0;
    assign rom[13'h0ec4] = 0;
    assign rom[13'h0ec5] = 0;
    assign rom[13'h0ec6] = 0;
    assign rom[13'h0ec7] = 0;
    assign rom[13'h0ec8] = 0;
    assign rom[13'h0ec9] = 0;
    assign rom[13'h0eca] = 0;
    assign rom[13'h0ecb] = 0;
    assign rom[13'h0ecc] = 0;
    assign rom[13'h0ecd] = 0;
    assign rom[13'h0ece] = 0;
    assign rom[13'h0ecf] = 0;
    assign rom[13'h0ed0] = 0;
    assign rom[13'h0ed1] = 0;
    assign rom[13'h0ed2] = 0;
    assign rom[13'h0ed3] = 1;
    assign rom[13'h0ed4] = 1;
    assign rom[13'h0ed5] = 0;
    assign rom[13'h0ed6] = 0;
    assign rom[13'h0ed7] = 0;
    assign rom[13'h0ed8] = 0;
    assign rom[13'h0ed9] = 0;
    assign rom[13'h0eda] = 0;
    assign rom[13'h0edb] = 1;
    assign rom[13'h0edc] = 1;
    assign rom[13'h0edd] = 0;
    assign rom[13'h0ede] = 0;
    assign rom[13'h0edf] = 0;
    assign rom[13'h0ee0] = 0;
    assign rom[13'h0ee1] = 0;
    assign rom[13'h0ee2] = 0;
    assign rom[13'h0ee3] = 0;
    assign rom[13'h0ee4] = 0;
    assign rom[13'h0ee5] = 0;
    assign rom[13'h0ee6] = 0;
    assign rom[13'h0ee7] = 0;
    assign rom[13'h0ee8] = 0;
    assign rom[13'h0ee9] = 0;
    assign rom[13'h0eea] = 0;
    assign rom[13'h0eeb] = 1;
    assign rom[13'h0eec] = 1;
    assign rom[13'h0eed] = 0;
    assign rom[13'h0eee] = 0;
    assign rom[13'h0eef] = 0;
    assign rom[13'h0ef0] = 0;
    assign rom[13'h0ef1] = 0;
    assign rom[13'h0ef2] = 0;
    assign rom[13'h0ef3] = 1;
    assign rom[13'h0ef4] = 1;
    assign rom[13'h0ef5] = 0;
    assign rom[13'h0ef6] = 0;
    assign rom[13'h0ef7] = 0;
    assign rom[13'h0ef8] = 0;
    assign rom[13'h0ef9] = 0;
    assign rom[13'h0efa] = 0;
    assign rom[13'h0efb] = 1;
    assign rom[13'h0efc] = 0;
    assign rom[13'h0efd] = 0;
    assign rom[13'h0efe] = 0;
    assign rom[13'h0eff] = 0;
    assign rom[13'h0f00] = 0;
    assign rom[13'h0f01] = 0;
    assign rom[13'h0f02] = 0;
    assign rom[13'h0f03] = 0;
    assign rom[13'h0f04] = 1;
    assign rom[13'h0f05] = 1;
    assign rom[13'h0f06] = 0;
    assign rom[13'h0f07] = 0;
    assign rom[13'h0f08] = 0;
    assign rom[13'h0f09] = 0;
    assign rom[13'h0f0a] = 0;
    assign rom[13'h0f0b] = 1;
    assign rom[13'h0f0c] = 1;
    assign rom[13'h0f0d] = 0;
    assign rom[13'h0f0e] = 0;
    assign rom[13'h0f0f] = 0;
    assign rom[13'h0f10] = 0;
    assign rom[13'h0f11] = 0;
    assign rom[13'h0f12] = 1;
    assign rom[13'h0f13] = 1;
    assign rom[13'h0f14] = 0;
    assign rom[13'h0f15] = 0;
    assign rom[13'h0f16] = 0;
    assign rom[13'h0f17] = 0;
    assign rom[13'h0f18] = 0;
    assign rom[13'h0f19] = 1;
    assign rom[13'h0f1a] = 1;
    assign rom[13'h0f1b] = 0;
    assign rom[13'h0f1c] = 0;
    assign rom[13'h0f1d] = 0;
    assign rom[13'h0f1e] = 0;
    assign rom[13'h0f1f] = 0;
    assign rom[13'h0f20] = 0;
    assign rom[13'h0f21] = 0;
    assign rom[13'h0f22] = 1;
    assign rom[13'h0f23] = 1;
    assign rom[13'h0f24] = 0;
    assign rom[13'h0f25] = 0;
    assign rom[13'h0f26] = 0;
    assign rom[13'h0f27] = 0;
    assign rom[13'h0f28] = 0;
    assign rom[13'h0f29] = 0;
    assign rom[13'h0f2a] = 0;
    assign rom[13'h0f2b] = 1;
    assign rom[13'h0f2c] = 1;
    assign rom[13'h0f2d] = 0;
    assign rom[13'h0f2e] = 0;
    assign rom[13'h0f2f] = 0;
    assign rom[13'h0f30] = 0;
    assign rom[13'h0f31] = 0;
    assign rom[13'h0f32] = 0;
    assign rom[13'h0f33] = 0;
    assign rom[13'h0f34] = 1;
    assign rom[13'h0f35] = 1;
    assign rom[13'h0f36] = 0;
    assign rom[13'h0f37] = 0;
    assign rom[13'h0f38] = 0;
    assign rom[13'h0f39] = 0;
    assign rom[13'h0f3a] = 0;
    assign rom[13'h0f3b] = 0;
    assign rom[13'h0f3c] = 0;
    assign rom[13'h0f3d] = 0;
    assign rom[13'h0f3e] = 0;
    assign rom[13'h0f3f] = 0;
    assign rom[13'h0f40] = 0;
    assign rom[13'h0f41] = 0;
    assign rom[13'h0f42] = 0;
    assign rom[13'h0f43] = 0;
    assign rom[13'h0f44] = 0;
    assign rom[13'h0f45] = 0;
    assign rom[13'h0f46] = 0;
    assign rom[13'h0f47] = 0;
    assign rom[13'h0f48] = 0;
    assign rom[13'h0f49] = 0;
    assign rom[13'h0f4a] = 0;
    assign rom[13'h0f4b] = 0;
    assign rom[13'h0f4c] = 0;
    assign rom[13'h0f4d] = 0;
    assign rom[13'h0f4e] = 0;
    assign rom[13'h0f4f] = 0;
    assign rom[13'h0f50] = 0;
    assign rom[13'h0f51] = 1;
    assign rom[13'h0f52] = 1;
    assign rom[13'h0f53] = 1;
    assign rom[13'h0f54] = 1;
    assign rom[13'h0f55] = 1;
    assign rom[13'h0f56] = 1;
    assign rom[13'h0f57] = 0;
    assign rom[13'h0f58] = 0;
    assign rom[13'h0f59] = 0;
    assign rom[13'h0f5a] = 0;
    assign rom[13'h0f5b] = 0;
    assign rom[13'h0f5c] = 0;
    assign rom[13'h0f5d] = 0;
    assign rom[13'h0f5e] = 0;
    assign rom[13'h0f5f] = 0;
    assign rom[13'h0f60] = 0;
    assign rom[13'h0f61] = 1;
    assign rom[13'h0f62] = 1;
    assign rom[13'h0f63] = 1;
    assign rom[13'h0f64] = 1;
    assign rom[13'h0f65] = 1;
    assign rom[13'h0f66] = 1;
    assign rom[13'h0f67] = 0;
    assign rom[13'h0f68] = 0;
    assign rom[13'h0f69] = 0;
    assign rom[13'h0f6a] = 0;
    assign rom[13'h0f6b] = 0;
    assign rom[13'h0f6c] = 0;
    assign rom[13'h0f6d] = 0;
    assign rom[13'h0f6e] = 0;
    assign rom[13'h0f6f] = 0;
    assign rom[13'h0f70] = 0;
    assign rom[13'h0f71] = 0;
    assign rom[13'h0f72] = 0;
    assign rom[13'h0f73] = 0;
    assign rom[13'h0f74] = 0;
    assign rom[13'h0f75] = 0;
    assign rom[13'h0f76] = 0;
    assign rom[13'h0f77] = 0;
    assign rom[13'h0f78] = 0;
    assign rom[13'h0f79] = 0;
    assign rom[13'h0f7a] = 0;
    assign rom[13'h0f7b] = 0;
    assign rom[13'h0f7c] = 0;
    assign rom[13'h0f7d] = 0;
    assign rom[13'h0f7e] = 0;
    assign rom[13'h0f7f] = 0;
    assign rom[13'h0f80] = 0;
    assign rom[13'h0f81] = 0;
    assign rom[13'h0f82] = 1;
    assign rom[13'h0f83] = 1;
    assign rom[13'h0f84] = 0;
    assign rom[13'h0f85] = 0;
    assign rom[13'h0f86] = 0;
    assign rom[13'h0f87] = 0;
    assign rom[13'h0f88] = 0;
    assign rom[13'h0f89] = 0;
    assign rom[13'h0f8a] = 0;
    assign rom[13'h0f8b] = 1;
    assign rom[13'h0f8c] = 1;
    assign rom[13'h0f8d] = 0;
    assign rom[13'h0f8e] = 0;
    assign rom[13'h0f8f] = 0;
    assign rom[13'h0f90] = 0;
    assign rom[13'h0f91] = 0;
    assign rom[13'h0f92] = 0;
    assign rom[13'h0f93] = 0;
    assign rom[13'h0f94] = 1;
    assign rom[13'h0f95] = 1;
    assign rom[13'h0f96] = 0;
    assign rom[13'h0f97] = 0;
    assign rom[13'h0f98] = 0;
    assign rom[13'h0f99] = 0;
    assign rom[13'h0f9a] = 0;
    assign rom[13'h0f9b] = 0;
    assign rom[13'h0f9c] = 0;
    assign rom[13'h0f9d] = 1;
    assign rom[13'h0f9e] = 1;
    assign rom[13'h0f9f] = 0;
    assign rom[13'h0fa0] = 0;
    assign rom[13'h0fa1] = 0;
    assign rom[13'h0fa2] = 0;
    assign rom[13'h0fa3] = 0;
    assign rom[13'h0fa4] = 1;
    assign rom[13'h0fa5] = 1;
    assign rom[13'h0fa6] = 0;
    assign rom[13'h0fa7] = 0;
    assign rom[13'h0fa8] = 0;
    assign rom[13'h0fa9] = 0;
    assign rom[13'h0faa] = 0;
    assign rom[13'h0fab] = 1;
    assign rom[13'h0fac] = 1;
    assign rom[13'h0fad] = 0;
    assign rom[13'h0fae] = 0;
    assign rom[13'h0faf] = 0;
    assign rom[13'h0fb0] = 0;
    assign rom[13'h0fb1] = 0;
    assign rom[13'h0fb2] = 1;
    assign rom[13'h0fb3] = 1;
    assign rom[13'h0fb4] = 0;
    assign rom[13'h0fb5] = 0;
    assign rom[13'h0fb6] = 0;
    assign rom[13'h0fb7] = 0;
    assign rom[13'h0fb8] = 0;
    assign rom[13'h0fb9] = 0;
    assign rom[13'h0fba] = 0;
    assign rom[13'h0fbb] = 0;
    assign rom[13'h0fbc] = 0;
    assign rom[13'h0fbd] = 0;
    assign rom[13'h0fbe] = 0;
    assign rom[13'h0fbf] = 0;
    assign rom[13'h0fc0] = 0;
    assign rom[13'h0fc1] = 0;
    assign rom[13'h0fc2] = 1;
    assign rom[13'h0fc3] = 1;
    assign rom[13'h0fc4] = 1;
    assign rom[13'h0fc5] = 1;
    assign rom[13'h0fc6] = 0;
    assign rom[13'h0fc7] = 0;
    assign rom[13'h0fc8] = 0;
    assign rom[13'h0fc9] = 1;
    assign rom[13'h0fca] = 1;
    assign rom[13'h0fcb] = 0;
    assign rom[13'h0fcc] = 0;
    assign rom[13'h0fcd] = 1;
    assign rom[13'h0fce] = 1;
    assign rom[13'h0fcf] = 0;
    assign rom[13'h0fd0] = 0;
    assign rom[13'h0fd1] = 0;
    assign rom[13'h0fd2] = 0;
    assign rom[13'h0fd3] = 0;
    assign rom[13'h0fd4] = 0;
    assign rom[13'h0fd5] = 1;
    assign rom[13'h0fd6] = 1;
    assign rom[13'h0fd7] = 0;
    assign rom[13'h0fd8] = 0;
    assign rom[13'h0fd9] = 0;
    assign rom[13'h0fda] = 0;
    assign rom[13'h0fdb] = 1;
    assign rom[13'h0fdc] = 1;
    assign rom[13'h0fdd] = 1;
    assign rom[13'h0fde] = 0;
    assign rom[13'h0fdf] = 0;
    assign rom[13'h0fe0] = 0;
    assign rom[13'h0fe1] = 0;
    assign rom[13'h0fe2] = 0;
    assign rom[13'h0fe3] = 1;
    assign rom[13'h0fe4] = 1;
    assign rom[13'h0fe5] = 0;
    assign rom[13'h0fe6] = 0;
    assign rom[13'h0fe7] = 0;
    assign rom[13'h0fe8] = 0;
    assign rom[13'h0fe9] = 0;
    assign rom[13'h0fea] = 0;
    assign rom[13'h0feb] = 0;
    assign rom[13'h0fec] = 0;
    assign rom[13'h0fed] = 0;
    assign rom[13'h0fee] = 0;
    assign rom[13'h0fef] = 0;
    assign rom[13'h0ff0] = 0;
    assign rom[13'h0ff1] = 0;
    assign rom[13'h0ff2] = 0;
    assign rom[13'h0ff3] = 1;
    assign rom[13'h0ff4] = 1;
    assign rom[13'h0ff5] = 0;
    assign rom[13'h0ff6] = 0;
    assign rom[13'h0ff7] = 0;
    assign rom[13'h0ff8] = 0;
    assign rom[13'h0ff9] = 0;
    assign rom[13'h0ffa] = 0;
    assign rom[13'h0ffb] = 0;
    assign rom[13'h0ffc] = 0;
    assign rom[13'h0ffd] = 0;
    assign rom[13'h0ffe] = 0;
    assign rom[13'h0fff] = 0;
    assign rom[13'h1000] = 0;
    assign rom[13'h1001] = 0;
    assign rom[13'h1002] = 1;
    assign rom[13'h1003] = 1;
    assign rom[13'h1004] = 1;
    assign rom[13'h1005] = 1;
    assign rom[13'h1006] = 0;
    assign rom[13'h1007] = 0;
    assign rom[13'h1008] = 0;
    assign rom[13'h1009] = 1;
    assign rom[13'h100a] = 1;
    assign rom[13'h100b] = 0;
    assign rom[13'h100c] = 0;
    assign rom[13'h100d] = 1;
    assign rom[13'h100e] = 1;
    assign rom[13'h100f] = 0;
    assign rom[13'h1010] = 0;
    assign rom[13'h1011] = 1;
    assign rom[13'h1012] = 1;
    assign rom[13'h1013] = 0;
    assign rom[13'h1014] = 1;
    assign rom[13'h1015] = 1;
    assign rom[13'h1016] = 1;
    assign rom[13'h1017] = 0;
    assign rom[13'h1018] = 0;
    assign rom[13'h1019] = 1;
    assign rom[13'h101a] = 1;
    assign rom[13'h101b] = 0;
    assign rom[13'h101c] = 1;
    assign rom[13'h101d] = 0;
    assign rom[13'h101e] = 1;
    assign rom[13'h101f] = 0;
    assign rom[13'h1020] = 0;
    assign rom[13'h1021] = 1;
    assign rom[13'h1022] = 1;
    assign rom[13'h1023] = 0;
    assign rom[13'h1024] = 1;
    assign rom[13'h1025] = 1;
    assign rom[13'h1026] = 1;
    assign rom[13'h1027] = 0;
    assign rom[13'h1028] = 0;
    assign rom[13'h1029] = 1;
    assign rom[13'h102a] = 1;
    assign rom[13'h102b] = 0;
    assign rom[13'h102c] = 0;
    assign rom[13'h102d] = 0;
    assign rom[13'h102e] = 0;
    assign rom[13'h102f] = 0;
    assign rom[13'h1030] = 0;
    assign rom[13'h1031] = 0;
    assign rom[13'h1032] = 1;
    assign rom[13'h1033] = 1;
    assign rom[13'h1034] = 1;
    assign rom[13'h1035] = 1;
    assign rom[13'h1036] = 1;
    assign rom[13'h1037] = 0;
    assign rom[13'h1038] = 0;
    assign rom[13'h1039] = 0;
    assign rom[13'h103a] = 0;
    assign rom[13'h103b] = 0;
    assign rom[13'h103c] = 0;
    assign rom[13'h103d] = 0;
    assign rom[13'h103e] = 0;
    assign rom[13'h103f] = 0;
    assign rom[13'h1040] = 0;
    assign rom[13'h1041] = 0;
    assign rom[13'h1042] = 1;
    assign rom[13'h1043] = 1;
    assign rom[13'h1044] = 1;
    assign rom[13'h1045] = 1;
    assign rom[13'h1046] = 0;
    assign rom[13'h1047] = 0;
    assign rom[13'h1048] = 0;
    assign rom[13'h1049] = 1;
    assign rom[13'h104a] = 1;
    assign rom[13'h104b] = 0;
    assign rom[13'h104c] = 0;
    assign rom[13'h104d] = 1;
    assign rom[13'h104e] = 1;
    assign rom[13'h104f] = 0;
    assign rom[13'h1050] = 0;
    assign rom[13'h1051] = 1;
    assign rom[13'h1052] = 1;
    assign rom[13'h1053] = 0;
    assign rom[13'h1054] = 0;
    assign rom[13'h1055] = 1;
    assign rom[13'h1056] = 1;
    assign rom[13'h1057] = 0;
    assign rom[13'h1058] = 0;
    assign rom[13'h1059] = 1;
    assign rom[13'h105a] = 1;
    assign rom[13'h105b] = 1;
    assign rom[13'h105c] = 1;
    assign rom[13'h105d] = 1;
    assign rom[13'h105e] = 1;
    assign rom[13'h105f] = 0;
    assign rom[13'h1060] = 0;
    assign rom[13'h1061] = 1;
    assign rom[13'h1062] = 1;
    assign rom[13'h1063] = 0;
    assign rom[13'h1064] = 0;
    assign rom[13'h1065] = 1;
    assign rom[13'h1066] = 1;
    assign rom[13'h1067] = 0;
    assign rom[13'h1068] = 0;
    assign rom[13'h1069] = 1;
    assign rom[13'h106a] = 1;
    assign rom[13'h106b] = 0;
    assign rom[13'h106c] = 0;
    assign rom[13'h106d] = 1;
    assign rom[13'h106e] = 1;
    assign rom[13'h106f] = 0;
    assign rom[13'h1070] = 0;
    assign rom[13'h1071] = 1;
    assign rom[13'h1072] = 1;
    assign rom[13'h1073] = 0;
    assign rom[13'h1074] = 0;
    assign rom[13'h1075] = 1;
    assign rom[13'h1076] = 1;
    assign rom[13'h1077] = 0;
    assign rom[13'h1078] = 0;
    assign rom[13'h1079] = 0;
    assign rom[13'h107a] = 0;
    assign rom[13'h107b] = 0;
    assign rom[13'h107c] = 0;
    assign rom[13'h107d] = 0;
    assign rom[13'h107e] = 0;
    assign rom[13'h107f] = 0;
    assign rom[13'h1080] = 0;
    assign rom[13'h1081] = 1;
    assign rom[13'h1082] = 1;
    assign rom[13'h1083] = 1;
    assign rom[13'h1084] = 1;
    assign rom[13'h1085] = 1;
    assign rom[13'h1086] = 0;
    assign rom[13'h1087] = 0;
    assign rom[13'h1088] = 0;
    assign rom[13'h1089] = 1;
    assign rom[13'h108a] = 1;
    assign rom[13'h108b] = 0;
    assign rom[13'h108c] = 0;
    assign rom[13'h108d] = 1;
    assign rom[13'h108e] = 1;
    assign rom[13'h108f] = 0;
    assign rom[13'h1090] = 0;
    assign rom[13'h1091] = 1;
    assign rom[13'h1092] = 1;
    assign rom[13'h1093] = 0;
    assign rom[13'h1094] = 0;
    assign rom[13'h1095] = 1;
    assign rom[13'h1096] = 1;
    assign rom[13'h1097] = 0;
    assign rom[13'h1098] = 0;
    assign rom[13'h1099] = 1;
    assign rom[13'h109a] = 1;
    assign rom[13'h109b] = 1;
    assign rom[13'h109c] = 1;
    assign rom[13'h109d] = 1;
    assign rom[13'h109e] = 0;
    assign rom[13'h109f] = 0;
    assign rom[13'h10a0] = 0;
    assign rom[13'h10a1] = 1;
    assign rom[13'h10a2] = 1;
    assign rom[13'h10a3] = 0;
    assign rom[13'h10a4] = 0;
    assign rom[13'h10a5] = 1;
    assign rom[13'h10a6] = 1;
    assign rom[13'h10a7] = 0;
    assign rom[13'h10a8] = 0;
    assign rom[13'h10a9] = 1;
    assign rom[13'h10aa] = 1;
    assign rom[13'h10ab] = 0;
    assign rom[13'h10ac] = 0;
    assign rom[13'h10ad] = 1;
    assign rom[13'h10ae] = 1;
    assign rom[13'h10af] = 0;
    assign rom[13'h10b0] = 0;
    assign rom[13'h10b1] = 1;
    assign rom[13'h10b2] = 1;
    assign rom[13'h10b3] = 1;
    assign rom[13'h10b4] = 1;
    assign rom[13'h10b5] = 1;
    assign rom[13'h10b6] = 0;
    assign rom[13'h10b7] = 0;
    assign rom[13'h10b8] = 0;
    assign rom[13'h10b9] = 0;
    assign rom[13'h10ba] = 0;
    assign rom[13'h10bb] = 0;
    assign rom[13'h10bc] = 0;
    assign rom[13'h10bd] = 0;
    assign rom[13'h10be] = 0;
    assign rom[13'h10bf] = 0;
    assign rom[13'h10c0] = 0;
    assign rom[13'h10c1] = 0;
    assign rom[13'h10c2] = 1;
    assign rom[13'h10c3] = 1;
    assign rom[13'h10c4] = 1;
    assign rom[13'h10c5] = 1;
    assign rom[13'h10c6] = 0;
    assign rom[13'h10c7] = 0;
    assign rom[13'h10c8] = 0;
    assign rom[13'h10c9] = 1;
    assign rom[13'h10ca] = 1;
    assign rom[13'h10cb] = 0;
    assign rom[13'h10cc] = 0;
    assign rom[13'h10cd] = 1;
    assign rom[13'h10ce] = 1;
    assign rom[13'h10cf] = 0;
    assign rom[13'h10d0] = 0;
    assign rom[13'h10d1] = 1;
    assign rom[13'h10d2] = 1;
    assign rom[13'h10d3] = 0;
    assign rom[13'h10d4] = 0;
    assign rom[13'h10d5] = 0;
    assign rom[13'h10d6] = 0;
    assign rom[13'h10d7] = 0;
    assign rom[13'h10d8] = 0;
    assign rom[13'h10d9] = 1;
    assign rom[13'h10da] = 1;
    assign rom[13'h10db] = 0;
    assign rom[13'h10dc] = 0;
    assign rom[13'h10dd] = 0;
    assign rom[13'h10de] = 0;
    assign rom[13'h10df] = 0;
    assign rom[13'h10e0] = 0;
    assign rom[13'h10e1] = 1;
    assign rom[13'h10e2] = 1;
    assign rom[13'h10e3] = 0;
    assign rom[13'h10e4] = 0;
    assign rom[13'h10e5] = 0;
    assign rom[13'h10e6] = 0;
    assign rom[13'h10e7] = 0;
    assign rom[13'h10e8] = 0;
    assign rom[13'h10e9] = 1;
    assign rom[13'h10ea] = 1;
    assign rom[13'h10eb] = 0;
    assign rom[13'h10ec] = 0;
    assign rom[13'h10ed] = 1;
    assign rom[13'h10ee] = 1;
    assign rom[13'h10ef] = 0;
    assign rom[13'h10f0] = 0;
    assign rom[13'h10f1] = 0;
    assign rom[13'h10f2] = 1;
    assign rom[13'h10f3] = 1;
    assign rom[13'h10f4] = 1;
    assign rom[13'h10f5] = 1;
    assign rom[13'h10f6] = 0;
    assign rom[13'h10f7] = 0;
    assign rom[13'h10f8] = 0;
    assign rom[13'h10f9] = 0;
    assign rom[13'h10fa] = 0;
    assign rom[13'h10fb] = 0;
    assign rom[13'h10fc] = 0;
    assign rom[13'h10fd] = 0;
    assign rom[13'h10fe] = 0;
    assign rom[13'h10ff] = 0;
    assign rom[13'h1100] = 0;
    assign rom[13'h1101] = 1;
    assign rom[13'h1102] = 1;
    assign rom[13'h1103] = 1;
    assign rom[13'h1104] = 1;
    assign rom[13'h1105] = 1;
    assign rom[13'h1106] = 0;
    assign rom[13'h1107] = 0;
    assign rom[13'h1108] = 0;
    assign rom[13'h1109] = 1;
    assign rom[13'h110a] = 1;
    assign rom[13'h110b] = 0;
    assign rom[13'h110c] = 0;
    assign rom[13'h110d] = 1;
    assign rom[13'h110e] = 1;
    assign rom[13'h110f] = 0;
    assign rom[13'h1110] = 0;
    assign rom[13'h1111] = 1;
    assign rom[13'h1112] = 1;
    assign rom[13'h1113] = 0;
    assign rom[13'h1114] = 0;
    assign rom[13'h1115] = 1;
    assign rom[13'h1116] = 1;
    assign rom[13'h1117] = 0;
    assign rom[13'h1118] = 0;
    assign rom[13'h1119] = 1;
    assign rom[13'h111a] = 1;
    assign rom[13'h111b] = 0;
    assign rom[13'h111c] = 0;
    assign rom[13'h111d] = 1;
    assign rom[13'h111e] = 1;
    assign rom[13'h111f] = 0;
    assign rom[13'h1120] = 0;
    assign rom[13'h1121] = 1;
    assign rom[13'h1122] = 1;
    assign rom[13'h1123] = 0;
    assign rom[13'h1124] = 0;
    assign rom[13'h1125] = 1;
    assign rom[13'h1126] = 1;
    assign rom[13'h1127] = 0;
    assign rom[13'h1128] = 0;
    assign rom[13'h1129] = 1;
    assign rom[13'h112a] = 1;
    assign rom[13'h112b] = 0;
    assign rom[13'h112c] = 0;
    assign rom[13'h112d] = 1;
    assign rom[13'h112e] = 1;
    assign rom[13'h112f] = 0;
    assign rom[13'h1130] = 0;
    assign rom[13'h1131] = 1;
    assign rom[13'h1132] = 1;
    assign rom[13'h1133] = 1;
    assign rom[13'h1134] = 1;
    assign rom[13'h1135] = 1;
    assign rom[13'h1136] = 0;
    assign rom[13'h1137] = 0;
    assign rom[13'h1138] = 0;
    assign rom[13'h1139] = 0;
    assign rom[13'h113a] = 0;
    assign rom[13'h113b] = 0;
    assign rom[13'h113c] = 0;
    assign rom[13'h113d] = 0;
    assign rom[13'h113e] = 0;
    assign rom[13'h113f] = 0;
    assign rom[13'h1140] = 0;
    assign rom[13'h1141] = 1;
    assign rom[13'h1142] = 1;
    assign rom[13'h1143] = 1;
    assign rom[13'h1144] = 1;
    assign rom[13'h1145] = 1;
    assign rom[13'h1146] = 1;
    assign rom[13'h1147] = 0;
    assign rom[13'h1148] = 0;
    assign rom[13'h1149] = 1;
    assign rom[13'h114a] = 1;
    assign rom[13'h114b] = 0;
    assign rom[13'h114c] = 0;
    assign rom[13'h114d] = 0;
    assign rom[13'h114e] = 0;
    assign rom[13'h114f] = 0;
    assign rom[13'h1150] = 0;
    assign rom[13'h1151] = 1;
    assign rom[13'h1152] = 1;
    assign rom[13'h1153] = 0;
    assign rom[13'h1154] = 0;
    assign rom[13'h1155] = 0;
    assign rom[13'h1156] = 0;
    assign rom[13'h1157] = 0;
    assign rom[13'h1158] = 0;
    assign rom[13'h1159] = 1;
    assign rom[13'h115a] = 1;
    assign rom[13'h115b] = 1;
    assign rom[13'h115c] = 1;
    assign rom[13'h115d] = 1;
    assign rom[13'h115e] = 0;
    assign rom[13'h115f] = 0;
    assign rom[13'h1160] = 0;
    assign rom[13'h1161] = 1;
    assign rom[13'h1162] = 1;
    assign rom[13'h1163] = 0;
    assign rom[13'h1164] = 0;
    assign rom[13'h1165] = 0;
    assign rom[13'h1166] = 0;
    assign rom[13'h1167] = 0;
    assign rom[13'h1168] = 0;
    assign rom[13'h1169] = 1;
    assign rom[13'h116a] = 1;
    assign rom[13'h116b] = 0;
    assign rom[13'h116c] = 0;
    assign rom[13'h116d] = 0;
    assign rom[13'h116e] = 0;
    assign rom[13'h116f] = 0;
    assign rom[13'h1170] = 0;
    assign rom[13'h1171] = 1;
    assign rom[13'h1172] = 1;
    assign rom[13'h1173] = 1;
    assign rom[13'h1174] = 1;
    assign rom[13'h1175] = 1;
    assign rom[13'h1176] = 1;
    assign rom[13'h1177] = 0;
    assign rom[13'h1178] = 0;
    assign rom[13'h1179] = 0;
    assign rom[13'h117a] = 0;
    assign rom[13'h117b] = 0;
    assign rom[13'h117c] = 0;
    assign rom[13'h117d] = 0;
    assign rom[13'h117e] = 0;
    assign rom[13'h117f] = 0;
    assign rom[13'h1180] = 0;
    assign rom[13'h1181] = 1;
    assign rom[13'h1182] = 1;
    assign rom[13'h1183] = 1;
    assign rom[13'h1184] = 1;
    assign rom[13'h1185] = 1;
    assign rom[13'h1186] = 1;
    assign rom[13'h1187] = 0;
    assign rom[13'h1188] = 0;
    assign rom[13'h1189] = 1;
    assign rom[13'h118a] = 1;
    assign rom[13'h118b] = 0;
    assign rom[13'h118c] = 0;
    assign rom[13'h118d] = 0;
    assign rom[13'h118e] = 0;
    assign rom[13'h118f] = 0;
    assign rom[13'h1190] = 0;
    assign rom[13'h1191] = 1;
    assign rom[13'h1192] = 1;
    assign rom[13'h1193] = 0;
    assign rom[13'h1194] = 0;
    assign rom[13'h1195] = 0;
    assign rom[13'h1196] = 0;
    assign rom[13'h1197] = 0;
    assign rom[13'h1198] = 0;
    assign rom[13'h1199] = 1;
    assign rom[13'h119a] = 1;
    assign rom[13'h119b] = 1;
    assign rom[13'h119c] = 1;
    assign rom[13'h119d] = 1;
    assign rom[13'h119e] = 0;
    assign rom[13'h119f] = 0;
    assign rom[13'h11a0] = 0;
    assign rom[13'h11a1] = 1;
    assign rom[13'h11a2] = 1;
    assign rom[13'h11a3] = 0;
    assign rom[13'h11a4] = 0;
    assign rom[13'h11a5] = 0;
    assign rom[13'h11a6] = 0;
    assign rom[13'h11a7] = 0;
    assign rom[13'h11a8] = 0;
    assign rom[13'h11a9] = 1;
    assign rom[13'h11aa] = 1;
    assign rom[13'h11ab] = 0;
    assign rom[13'h11ac] = 0;
    assign rom[13'h11ad] = 0;
    assign rom[13'h11ae] = 0;
    assign rom[13'h11af] = 0;
    assign rom[13'h11b0] = 0;
    assign rom[13'h11b1] = 1;
    assign rom[13'h11b2] = 1;
    assign rom[13'h11b3] = 0;
    assign rom[13'h11b4] = 0;
    assign rom[13'h11b5] = 0;
    assign rom[13'h11b6] = 0;
    assign rom[13'h11b7] = 0;
    assign rom[13'h11b8] = 0;
    assign rom[13'h11b9] = 0;
    assign rom[13'h11ba] = 0;
    assign rom[13'h11bb] = 0;
    assign rom[13'h11bc] = 0;
    assign rom[13'h11bd] = 0;
    assign rom[13'h11be] = 0;
    assign rom[13'h11bf] = 0;
    assign rom[13'h11c0] = 0;
    assign rom[13'h11c1] = 0;
    assign rom[13'h11c2] = 1;
    assign rom[13'h11c3] = 1;
    assign rom[13'h11c4] = 1;
    assign rom[13'h11c5] = 1;
    assign rom[13'h11c6] = 0;
    assign rom[13'h11c7] = 0;
    assign rom[13'h11c8] = 0;
    assign rom[13'h11c9] = 1;
    assign rom[13'h11ca] = 1;
    assign rom[13'h11cb] = 0;
    assign rom[13'h11cc] = 0;
    assign rom[13'h11cd] = 1;
    assign rom[13'h11ce] = 1;
    assign rom[13'h11cf] = 0;
    assign rom[13'h11d0] = 0;
    assign rom[13'h11d1] = 1;
    assign rom[13'h11d2] = 1;
    assign rom[13'h11d3] = 0;
    assign rom[13'h11d4] = 0;
    assign rom[13'h11d5] = 0;
    assign rom[13'h11d6] = 0;
    assign rom[13'h11d7] = 0;
    assign rom[13'h11d8] = 0;
    assign rom[13'h11d9] = 1;
    assign rom[13'h11da] = 1;
    assign rom[13'h11db] = 0;
    assign rom[13'h11dc] = 1;
    assign rom[13'h11dd] = 1;
    assign rom[13'h11de] = 1;
    assign rom[13'h11df] = 0;
    assign rom[13'h11e0] = 0;
    assign rom[13'h11e1] = 1;
    assign rom[13'h11e2] = 1;
    assign rom[13'h11e3] = 0;
    assign rom[13'h11e4] = 0;
    assign rom[13'h11e5] = 1;
    assign rom[13'h11e6] = 1;
    assign rom[13'h11e7] = 0;
    assign rom[13'h11e8] = 0;
    assign rom[13'h11e9] = 1;
    assign rom[13'h11ea] = 1;
    assign rom[13'h11eb] = 0;
    assign rom[13'h11ec] = 0;
    assign rom[13'h11ed] = 1;
    assign rom[13'h11ee] = 1;
    assign rom[13'h11ef] = 0;
    assign rom[13'h11f0] = 0;
    assign rom[13'h11f1] = 0;
    assign rom[13'h11f2] = 1;
    assign rom[13'h11f3] = 1;
    assign rom[13'h11f4] = 1;
    assign rom[13'h11f5] = 1;
    assign rom[13'h11f6] = 0;
    assign rom[13'h11f7] = 0;
    assign rom[13'h11f8] = 0;
    assign rom[13'h11f9] = 0;
    assign rom[13'h11fa] = 0;
    assign rom[13'h11fb] = 0;
    assign rom[13'h11fc] = 0;
    assign rom[13'h11fd] = 0;
    assign rom[13'h11fe] = 0;
    assign rom[13'h11ff] = 0;
    assign rom[13'h1200] = 0;
    assign rom[13'h1201] = 1;
    assign rom[13'h1202] = 1;
    assign rom[13'h1203] = 0;
    assign rom[13'h1204] = 0;
    assign rom[13'h1205] = 1;
    assign rom[13'h1206] = 1;
    assign rom[13'h1207] = 0;
    assign rom[13'h1208] = 0;
    assign rom[13'h1209] = 1;
    assign rom[13'h120a] = 1;
    assign rom[13'h120b] = 0;
    assign rom[13'h120c] = 0;
    assign rom[13'h120d] = 1;
    assign rom[13'h120e] = 1;
    assign rom[13'h120f] = 0;
    assign rom[13'h1210] = 0;
    assign rom[13'h1211] = 1;
    assign rom[13'h1212] = 1;
    assign rom[13'h1213] = 0;
    assign rom[13'h1214] = 0;
    assign rom[13'h1215] = 1;
    assign rom[13'h1216] = 1;
    assign rom[13'h1217] = 0;
    assign rom[13'h1218] = 0;
    assign rom[13'h1219] = 1;
    assign rom[13'h121a] = 1;
    assign rom[13'h121b] = 1;
    assign rom[13'h121c] = 1;
    assign rom[13'h121d] = 1;
    assign rom[13'h121e] = 1;
    assign rom[13'h121f] = 0;
    assign rom[13'h1220] = 0;
    assign rom[13'h1221] = 1;
    assign rom[13'h1222] = 1;
    assign rom[13'h1223] = 0;
    assign rom[13'h1224] = 0;
    assign rom[13'h1225] = 1;
    assign rom[13'h1226] = 1;
    assign rom[13'h1227] = 0;
    assign rom[13'h1228] = 0;
    assign rom[13'h1229] = 1;
    assign rom[13'h122a] = 1;
    assign rom[13'h122b] = 0;
    assign rom[13'h122c] = 0;
    assign rom[13'h122d] = 1;
    assign rom[13'h122e] = 1;
    assign rom[13'h122f] = 0;
    assign rom[13'h1230] = 0;
    assign rom[13'h1231] = 1;
    assign rom[13'h1232] = 1;
    assign rom[13'h1233] = 0;
    assign rom[13'h1234] = 0;
    assign rom[13'h1235] = 1;
    assign rom[13'h1236] = 1;
    assign rom[13'h1237] = 0;
    assign rom[13'h1238] = 0;
    assign rom[13'h1239] = 0;
    assign rom[13'h123a] = 0;
    assign rom[13'h123b] = 0;
    assign rom[13'h123c] = 0;
    assign rom[13'h123d] = 0;
    assign rom[13'h123e] = 0;
    assign rom[13'h123f] = 0;
    assign rom[13'h1240] = 0;
    assign rom[13'h1241] = 0;
    assign rom[13'h1242] = 1;
    assign rom[13'h1243] = 1;
    assign rom[13'h1244] = 1;
    assign rom[13'h1245] = 1;
    assign rom[13'h1246] = 0;
    assign rom[13'h1247] = 0;
    assign rom[13'h1248] = 0;
    assign rom[13'h1249] = 0;
    assign rom[13'h124a] = 0;
    assign rom[13'h124b] = 1;
    assign rom[13'h124c] = 1;
    assign rom[13'h124d] = 0;
    assign rom[13'h124e] = 0;
    assign rom[13'h124f] = 0;
    assign rom[13'h1250] = 0;
    assign rom[13'h1251] = 0;
    assign rom[13'h1252] = 0;
    assign rom[13'h1253] = 1;
    assign rom[13'h1254] = 1;
    assign rom[13'h1255] = 0;
    assign rom[13'h1256] = 0;
    assign rom[13'h1257] = 0;
    assign rom[13'h1258] = 0;
    assign rom[13'h1259] = 0;
    assign rom[13'h125a] = 0;
    assign rom[13'h125b] = 1;
    assign rom[13'h125c] = 1;
    assign rom[13'h125d] = 0;
    assign rom[13'h125e] = 0;
    assign rom[13'h125f] = 0;
    assign rom[13'h1260] = 0;
    assign rom[13'h1261] = 0;
    assign rom[13'h1262] = 0;
    assign rom[13'h1263] = 1;
    assign rom[13'h1264] = 1;
    assign rom[13'h1265] = 0;
    assign rom[13'h1266] = 0;
    assign rom[13'h1267] = 0;
    assign rom[13'h1268] = 0;
    assign rom[13'h1269] = 0;
    assign rom[13'h126a] = 0;
    assign rom[13'h126b] = 1;
    assign rom[13'h126c] = 1;
    assign rom[13'h126d] = 0;
    assign rom[13'h126e] = 0;
    assign rom[13'h126f] = 0;
    assign rom[13'h1270] = 0;
    assign rom[13'h1271] = 0;
    assign rom[13'h1272] = 1;
    assign rom[13'h1273] = 1;
    assign rom[13'h1274] = 1;
    assign rom[13'h1275] = 1;
    assign rom[13'h1276] = 0;
    assign rom[13'h1277] = 0;
    assign rom[13'h1278] = 0;
    assign rom[13'h1279] = 0;
    assign rom[13'h127a] = 0;
    assign rom[13'h127b] = 0;
    assign rom[13'h127c] = 0;
    assign rom[13'h127d] = 0;
    assign rom[13'h127e] = 0;
    assign rom[13'h127f] = 0;
    assign rom[13'h1280] = 0;
    assign rom[13'h1281] = 0;
    assign rom[13'h1282] = 1;
    assign rom[13'h1283] = 1;
    assign rom[13'h1284] = 1;
    assign rom[13'h1285] = 1;
    assign rom[13'h1286] = 1;
    assign rom[13'h1287] = 0;
    assign rom[13'h1288] = 0;
    assign rom[13'h1289] = 0;
    assign rom[13'h128a] = 0;
    assign rom[13'h128b] = 0;
    assign rom[13'h128c] = 1;
    assign rom[13'h128d] = 1;
    assign rom[13'h128e] = 0;
    assign rom[13'h128f] = 0;
    assign rom[13'h1290] = 0;
    assign rom[13'h1291] = 0;
    assign rom[13'h1292] = 0;
    assign rom[13'h1293] = 0;
    assign rom[13'h1294] = 1;
    assign rom[13'h1295] = 1;
    assign rom[13'h1296] = 0;
    assign rom[13'h1297] = 0;
    assign rom[13'h1298] = 0;
    assign rom[13'h1299] = 0;
    assign rom[13'h129a] = 0;
    assign rom[13'h129b] = 0;
    assign rom[13'h129c] = 1;
    assign rom[13'h129d] = 1;
    assign rom[13'h129e] = 0;
    assign rom[13'h129f] = 0;
    assign rom[13'h12a0] = 0;
    assign rom[13'h12a1] = 0;
    assign rom[13'h12a2] = 0;
    assign rom[13'h12a3] = 0;
    assign rom[13'h12a4] = 1;
    assign rom[13'h12a5] = 1;
    assign rom[13'h12a6] = 0;
    assign rom[13'h12a7] = 0;
    assign rom[13'h12a8] = 0;
    assign rom[13'h12a9] = 1;
    assign rom[13'h12aa] = 1;
    assign rom[13'h12ab] = 0;
    assign rom[13'h12ac] = 1;
    assign rom[13'h12ad] = 1;
    assign rom[13'h12ae] = 0;
    assign rom[13'h12af] = 0;
    assign rom[13'h12b0] = 0;
    assign rom[13'h12b1] = 0;
    assign rom[13'h12b2] = 1;
    assign rom[13'h12b3] = 1;
    assign rom[13'h12b4] = 1;
    assign rom[13'h12b5] = 0;
    assign rom[13'h12b6] = 0;
    assign rom[13'h12b7] = 0;
    assign rom[13'h12b8] = 0;
    assign rom[13'h12b9] = 0;
    assign rom[13'h12ba] = 0;
    assign rom[13'h12bb] = 0;
    assign rom[13'h12bc] = 0;
    assign rom[13'h12bd] = 0;
    assign rom[13'h12be] = 0;
    assign rom[13'h12bf] = 0;
    assign rom[13'h12c0] = 0;
    assign rom[13'h12c1] = 1;
    assign rom[13'h12c2] = 1;
    assign rom[13'h12c3] = 0;
    assign rom[13'h12c4] = 0;
    assign rom[13'h12c5] = 1;
    assign rom[13'h12c6] = 1;
    assign rom[13'h12c7] = 0;
    assign rom[13'h12c8] = 0;
    assign rom[13'h12c9] = 1;
    assign rom[13'h12ca] = 1;
    assign rom[13'h12cb] = 0;
    assign rom[13'h12cc] = 1;
    assign rom[13'h12cd] = 1;
    assign rom[13'h12ce] = 0;
    assign rom[13'h12cf] = 0;
    assign rom[13'h12d0] = 0;
    assign rom[13'h12d1] = 1;
    assign rom[13'h12d2] = 1;
    assign rom[13'h12d3] = 1;
    assign rom[13'h12d4] = 1;
    assign rom[13'h12d5] = 0;
    assign rom[13'h12d6] = 0;
    assign rom[13'h12d7] = 0;
    assign rom[13'h12d8] = 0;
    assign rom[13'h12d9] = 1;
    assign rom[13'h12da] = 1;
    assign rom[13'h12db] = 1;
    assign rom[13'h12dc] = 0;
    assign rom[13'h12dd] = 0;
    assign rom[13'h12de] = 0;
    assign rom[13'h12df] = 0;
    assign rom[13'h12e0] = 0;
    assign rom[13'h12e1] = 1;
    assign rom[13'h12e2] = 1;
    assign rom[13'h12e3] = 1;
    assign rom[13'h12e4] = 1;
    assign rom[13'h12e5] = 0;
    assign rom[13'h12e6] = 0;
    assign rom[13'h12e7] = 0;
    assign rom[13'h12e8] = 0;
    assign rom[13'h12e9] = 1;
    assign rom[13'h12ea] = 1;
    assign rom[13'h12eb] = 0;
    assign rom[13'h12ec] = 1;
    assign rom[13'h12ed] = 1;
    assign rom[13'h12ee] = 0;
    assign rom[13'h12ef] = 0;
    assign rom[13'h12f0] = 0;
    assign rom[13'h12f1] = 1;
    assign rom[13'h12f2] = 1;
    assign rom[13'h12f3] = 0;
    assign rom[13'h12f4] = 0;
    assign rom[13'h12f5] = 1;
    assign rom[13'h12f6] = 1;
    assign rom[13'h12f7] = 0;
    assign rom[13'h12f8] = 0;
    assign rom[13'h12f9] = 0;
    assign rom[13'h12fa] = 0;
    assign rom[13'h12fb] = 0;
    assign rom[13'h12fc] = 0;
    assign rom[13'h12fd] = 0;
    assign rom[13'h12fe] = 0;
    assign rom[13'h12ff] = 0;
    assign rom[13'h1300] = 0;
    assign rom[13'h1301] = 1;
    assign rom[13'h1302] = 1;
    assign rom[13'h1303] = 0;
    assign rom[13'h1304] = 0;
    assign rom[13'h1305] = 0;
    assign rom[13'h1306] = 0;
    assign rom[13'h1307] = 0;
    assign rom[13'h1308] = 0;
    assign rom[13'h1309] = 1;
    assign rom[13'h130a] = 1;
    assign rom[13'h130b] = 0;
    assign rom[13'h130c] = 0;
    assign rom[13'h130d] = 0;
    assign rom[13'h130e] = 0;
    assign rom[13'h130f] = 0;
    assign rom[13'h1310] = 0;
    assign rom[13'h1311] = 1;
    assign rom[13'h1312] = 1;
    assign rom[13'h1313] = 0;
    assign rom[13'h1314] = 0;
    assign rom[13'h1315] = 0;
    assign rom[13'h1316] = 0;
    assign rom[13'h1317] = 0;
    assign rom[13'h1318] = 0;
    assign rom[13'h1319] = 1;
    assign rom[13'h131a] = 1;
    assign rom[13'h131b] = 0;
    assign rom[13'h131c] = 0;
    assign rom[13'h131d] = 0;
    assign rom[13'h131e] = 0;
    assign rom[13'h131f] = 0;
    assign rom[13'h1320] = 0;
    assign rom[13'h1321] = 1;
    assign rom[13'h1322] = 1;
    assign rom[13'h1323] = 0;
    assign rom[13'h1324] = 0;
    assign rom[13'h1325] = 0;
    assign rom[13'h1326] = 0;
    assign rom[13'h1327] = 0;
    assign rom[13'h1328] = 0;
    assign rom[13'h1329] = 1;
    assign rom[13'h132a] = 1;
    assign rom[13'h132b] = 0;
    assign rom[13'h132c] = 0;
    assign rom[13'h132d] = 0;
    assign rom[13'h132e] = 0;
    assign rom[13'h132f] = 0;
    assign rom[13'h1330] = 0;
    assign rom[13'h1331] = 1;
    assign rom[13'h1332] = 1;
    assign rom[13'h1333] = 1;
    assign rom[13'h1334] = 1;
    assign rom[13'h1335] = 1;
    assign rom[13'h1336] = 1;
    assign rom[13'h1337] = 0;
    assign rom[13'h1338] = 0;
    assign rom[13'h1339] = 0;
    assign rom[13'h133a] = 0;
    assign rom[13'h133b] = 0;
    assign rom[13'h133c] = 0;
    assign rom[13'h133d] = 0;
    assign rom[13'h133e] = 0;
    assign rom[13'h133f] = 0;
    assign rom[13'h1340] = 1;
    assign rom[13'h1341] = 1;
    assign rom[13'h1342] = 0;
    assign rom[13'h1343] = 0;
    assign rom[13'h1344] = 0;
    assign rom[13'h1345] = 1;
    assign rom[13'h1346] = 1;
    assign rom[13'h1347] = 0;
    assign rom[13'h1348] = 1;
    assign rom[13'h1349] = 1;
    assign rom[13'h134a] = 1;
    assign rom[13'h134b] = 0;
    assign rom[13'h134c] = 1;
    assign rom[13'h134d] = 1;
    assign rom[13'h134e] = 1;
    assign rom[13'h134f] = 0;
    assign rom[13'h1350] = 1;
    assign rom[13'h1351] = 1;
    assign rom[13'h1352] = 1;
    assign rom[13'h1353] = 1;
    assign rom[13'h1354] = 1;
    assign rom[13'h1355] = 1;
    assign rom[13'h1356] = 1;
    assign rom[13'h1357] = 0;
    assign rom[13'h1358] = 1;
    assign rom[13'h1359] = 1;
    assign rom[13'h135a] = 0;
    assign rom[13'h135b] = 1;
    assign rom[13'h135c] = 0;
    assign rom[13'h135d] = 1;
    assign rom[13'h135e] = 1;
    assign rom[13'h135f] = 0;
    assign rom[13'h1360] = 1;
    assign rom[13'h1361] = 1;
    assign rom[13'h1362] = 0;
    assign rom[13'h1363] = 0;
    assign rom[13'h1364] = 0;
    assign rom[13'h1365] = 1;
    assign rom[13'h1366] = 1;
    assign rom[13'h1367] = 0;
    assign rom[13'h1368] = 1;
    assign rom[13'h1369] = 1;
    assign rom[13'h136a] = 0;
    assign rom[13'h136b] = 0;
    assign rom[13'h136c] = 0;
    assign rom[13'h136d] = 1;
    assign rom[13'h136e] = 1;
    assign rom[13'h136f] = 0;
    assign rom[13'h1370] = 1;
    assign rom[13'h1371] = 1;
    assign rom[13'h1372] = 0;
    assign rom[13'h1373] = 0;
    assign rom[13'h1374] = 0;
    assign rom[13'h1375] = 1;
    assign rom[13'h1376] = 1;
    assign rom[13'h1377] = 0;
    assign rom[13'h1378] = 0;
    assign rom[13'h1379] = 0;
    assign rom[13'h137a] = 0;
    assign rom[13'h137b] = 0;
    assign rom[13'h137c] = 0;
    assign rom[13'h137d] = 0;
    assign rom[13'h137e] = 0;
    assign rom[13'h137f] = 0;
    assign rom[13'h1380] = 0;
    assign rom[13'h1381] = 1;
    assign rom[13'h1382] = 1;
    assign rom[13'h1383] = 0;
    assign rom[13'h1384] = 0;
    assign rom[13'h1385] = 1;
    assign rom[13'h1386] = 1;
    assign rom[13'h1387] = 0;
    assign rom[13'h1388] = 0;
    assign rom[13'h1389] = 1;
    assign rom[13'h138a] = 1;
    assign rom[13'h138b] = 0;
    assign rom[13'h138c] = 0;
    assign rom[13'h138d] = 1;
    assign rom[13'h138e] = 1;
    assign rom[13'h138f] = 0;
    assign rom[13'h1390] = 0;
    assign rom[13'h1391] = 1;
    assign rom[13'h1392] = 1;
    assign rom[13'h1393] = 1;
    assign rom[13'h1394] = 0;
    assign rom[13'h1395] = 1;
    assign rom[13'h1396] = 1;
    assign rom[13'h1397] = 0;
    assign rom[13'h1398] = 0;
    assign rom[13'h1399] = 1;
    assign rom[13'h139a] = 1;
    assign rom[13'h139b] = 1;
    assign rom[13'h139c] = 1;
    assign rom[13'h139d] = 1;
    assign rom[13'h139e] = 1;
    assign rom[13'h139f] = 0;
    assign rom[13'h13a0] = 0;
    assign rom[13'h13a1] = 1;
    assign rom[13'h13a2] = 1;
    assign rom[13'h13a3] = 0;
    assign rom[13'h13a4] = 1;
    assign rom[13'h13a5] = 1;
    assign rom[13'h13a6] = 1;
    assign rom[13'h13a7] = 0;
    assign rom[13'h13a8] = 0;
    assign rom[13'h13a9] = 1;
    assign rom[13'h13aa] = 1;
    assign rom[13'h13ab] = 0;
    assign rom[13'h13ac] = 0;
    assign rom[13'h13ad] = 1;
    assign rom[13'h13ae] = 1;
    assign rom[13'h13af] = 0;
    assign rom[13'h13b0] = 0;
    assign rom[13'h13b1] = 1;
    assign rom[13'h13b2] = 1;
    assign rom[13'h13b3] = 0;
    assign rom[13'h13b4] = 0;
    assign rom[13'h13b5] = 1;
    assign rom[13'h13b6] = 1;
    assign rom[13'h13b7] = 0;
    assign rom[13'h13b8] = 0;
    assign rom[13'h13b9] = 0;
    assign rom[13'h13ba] = 0;
    assign rom[13'h13bb] = 0;
    assign rom[13'h13bc] = 0;
    assign rom[13'h13bd] = 0;
    assign rom[13'h13be] = 0;
    assign rom[13'h13bf] = 0;
    assign rom[13'h13c0] = 0;
    assign rom[13'h13c1] = 0;
    assign rom[13'h13c2] = 1;
    assign rom[13'h13c3] = 1;
    assign rom[13'h13c4] = 1;
    assign rom[13'h13c5] = 1;
    assign rom[13'h13c6] = 0;
    assign rom[13'h13c7] = 0;
    assign rom[13'h13c8] = 0;
    assign rom[13'h13c9] = 1;
    assign rom[13'h13ca] = 1;
    assign rom[13'h13cb] = 0;
    assign rom[13'h13cc] = 0;
    assign rom[13'h13cd] = 1;
    assign rom[13'h13ce] = 1;
    assign rom[13'h13cf] = 0;
    assign rom[13'h13d0] = 0;
    assign rom[13'h13d1] = 1;
    assign rom[13'h13d2] = 1;
    assign rom[13'h13d3] = 0;
    assign rom[13'h13d4] = 0;
    assign rom[13'h13d5] = 1;
    assign rom[13'h13d6] = 1;
    assign rom[13'h13d7] = 0;
    assign rom[13'h13d8] = 0;
    assign rom[13'h13d9] = 1;
    assign rom[13'h13da] = 1;
    assign rom[13'h13db] = 0;
    assign rom[13'h13dc] = 0;
    assign rom[13'h13dd] = 1;
    assign rom[13'h13de] = 1;
    assign rom[13'h13df] = 0;
    assign rom[13'h13e0] = 0;
    assign rom[13'h13e1] = 1;
    assign rom[13'h13e2] = 1;
    assign rom[13'h13e3] = 0;
    assign rom[13'h13e4] = 0;
    assign rom[13'h13e5] = 1;
    assign rom[13'h13e6] = 1;
    assign rom[13'h13e7] = 0;
    assign rom[13'h13e8] = 0;
    assign rom[13'h13e9] = 1;
    assign rom[13'h13ea] = 1;
    assign rom[13'h13eb] = 0;
    assign rom[13'h13ec] = 0;
    assign rom[13'h13ed] = 1;
    assign rom[13'h13ee] = 1;
    assign rom[13'h13ef] = 0;
    assign rom[13'h13f0] = 0;
    assign rom[13'h13f1] = 0;
    assign rom[13'h13f2] = 1;
    assign rom[13'h13f3] = 1;
    assign rom[13'h13f4] = 1;
    assign rom[13'h13f5] = 1;
    assign rom[13'h13f6] = 0;
    assign rom[13'h13f7] = 0;
    assign rom[13'h13f8] = 0;
    assign rom[13'h13f9] = 0;
    assign rom[13'h13fa] = 0;
    assign rom[13'h13fb] = 0;
    assign rom[13'h13fc] = 0;
    assign rom[13'h13fd] = 0;
    assign rom[13'h13fe] = 0;
    assign rom[13'h13ff] = 0;
    assign rom[13'h1400] = 0;
    assign rom[13'h1401] = 1;
    assign rom[13'h1402] = 1;
    assign rom[13'h1403] = 1;
    assign rom[13'h1404] = 1;
    assign rom[13'h1405] = 1;
    assign rom[13'h1406] = 0;
    assign rom[13'h1407] = 0;
    assign rom[13'h1408] = 0;
    assign rom[13'h1409] = 1;
    assign rom[13'h140a] = 1;
    assign rom[13'h140b] = 0;
    assign rom[13'h140c] = 0;
    assign rom[13'h140d] = 1;
    assign rom[13'h140e] = 1;
    assign rom[13'h140f] = 0;
    assign rom[13'h1410] = 0;
    assign rom[13'h1411] = 1;
    assign rom[13'h1412] = 1;
    assign rom[13'h1413] = 0;
    assign rom[13'h1414] = 0;
    assign rom[13'h1415] = 1;
    assign rom[13'h1416] = 1;
    assign rom[13'h1417] = 0;
    assign rom[13'h1418] = 0;
    assign rom[13'h1419] = 1;
    assign rom[13'h141a] = 1;
    assign rom[13'h141b] = 1;
    assign rom[13'h141c] = 1;
    assign rom[13'h141d] = 1;
    assign rom[13'h141e] = 0;
    assign rom[13'h141f] = 0;
    assign rom[13'h1420] = 0;
    assign rom[13'h1421] = 1;
    assign rom[13'h1422] = 1;
    assign rom[13'h1423] = 0;
    assign rom[13'h1424] = 0;
    assign rom[13'h1425] = 0;
    assign rom[13'h1426] = 0;
    assign rom[13'h1427] = 0;
    assign rom[13'h1428] = 0;
    assign rom[13'h1429] = 1;
    assign rom[13'h142a] = 1;
    assign rom[13'h142b] = 0;
    assign rom[13'h142c] = 0;
    assign rom[13'h142d] = 0;
    assign rom[13'h142e] = 0;
    assign rom[13'h142f] = 0;
    assign rom[13'h1430] = 0;
    assign rom[13'h1431] = 1;
    assign rom[13'h1432] = 1;
    assign rom[13'h1433] = 0;
    assign rom[13'h1434] = 0;
    assign rom[13'h1435] = 0;
    assign rom[13'h1436] = 0;
    assign rom[13'h1437] = 0;
    assign rom[13'h1438] = 0;
    assign rom[13'h1439] = 0;
    assign rom[13'h143a] = 0;
    assign rom[13'h143b] = 0;
    assign rom[13'h143c] = 0;
    assign rom[13'h143d] = 0;
    assign rom[13'h143e] = 0;
    assign rom[13'h143f] = 0;
    assign rom[13'h1440] = 0;
    assign rom[13'h1441] = 0;
    assign rom[13'h1442] = 1;
    assign rom[13'h1443] = 1;
    assign rom[13'h1444] = 1;
    assign rom[13'h1445] = 1;
    assign rom[13'h1446] = 0;
    assign rom[13'h1447] = 0;
    assign rom[13'h1448] = 0;
    assign rom[13'h1449] = 1;
    assign rom[13'h144a] = 1;
    assign rom[13'h144b] = 0;
    assign rom[13'h144c] = 0;
    assign rom[13'h144d] = 1;
    assign rom[13'h144e] = 1;
    assign rom[13'h144f] = 0;
    assign rom[13'h1450] = 0;
    assign rom[13'h1451] = 1;
    assign rom[13'h1452] = 1;
    assign rom[13'h1453] = 0;
    assign rom[13'h1454] = 0;
    assign rom[13'h1455] = 1;
    assign rom[13'h1456] = 1;
    assign rom[13'h1457] = 0;
    assign rom[13'h1458] = 0;
    assign rom[13'h1459] = 1;
    assign rom[13'h145a] = 1;
    assign rom[13'h145b] = 0;
    assign rom[13'h145c] = 0;
    assign rom[13'h145d] = 1;
    assign rom[13'h145e] = 1;
    assign rom[13'h145f] = 0;
    assign rom[13'h1460] = 0;
    assign rom[13'h1461] = 1;
    assign rom[13'h1462] = 1;
    assign rom[13'h1463] = 0;
    assign rom[13'h1464] = 1;
    assign rom[13'h1465] = 1;
    assign rom[13'h1466] = 1;
    assign rom[13'h1467] = 0;
    assign rom[13'h1468] = 0;
    assign rom[13'h1469] = 1;
    assign rom[13'h146a] = 1;
    assign rom[13'h146b] = 0;
    assign rom[13'h146c] = 0;
    assign rom[13'h146d] = 1;
    assign rom[13'h146e] = 1;
    assign rom[13'h146f] = 0;
    assign rom[13'h1470] = 0;
    assign rom[13'h1471] = 0;
    assign rom[13'h1472] = 1;
    assign rom[13'h1473] = 1;
    assign rom[13'h1474] = 1;
    assign rom[13'h1475] = 1;
    assign rom[13'h1476] = 1;
    assign rom[13'h1477] = 0;
    assign rom[13'h1478] = 0;
    assign rom[13'h1479] = 0;
    assign rom[13'h147a] = 0;
    assign rom[13'h147b] = 0;
    assign rom[13'h147c] = 0;
    assign rom[13'h147d] = 0;
    assign rom[13'h147e] = 0;
    assign rom[13'h147f] = 0;
    assign rom[13'h1480] = 0;
    assign rom[13'h1481] = 1;
    assign rom[13'h1482] = 1;
    assign rom[13'h1483] = 1;
    assign rom[13'h1484] = 1;
    assign rom[13'h1485] = 1;
    assign rom[13'h1486] = 0;
    assign rom[13'h1487] = 0;
    assign rom[13'h1488] = 0;
    assign rom[13'h1489] = 1;
    assign rom[13'h148a] = 1;
    assign rom[13'h148b] = 0;
    assign rom[13'h148c] = 0;
    assign rom[13'h148d] = 1;
    assign rom[13'h148e] = 1;
    assign rom[13'h148f] = 0;
    assign rom[13'h1490] = 0;
    assign rom[13'h1491] = 1;
    assign rom[13'h1492] = 1;
    assign rom[13'h1493] = 0;
    assign rom[13'h1494] = 0;
    assign rom[13'h1495] = 1;
    assign rom[13'h1496] = 1;
    assign rom[13'h1497] = 0;
    assign rom[13'h1498] = 0;
    assign rom[13'h1499] = 1;
    assign rom[13'h149a] = 1;
    assign rom[13'h149b] = 1;
    assign rom[13'h149c] = 1;
    assign rom[13'h149d] = 1;
    assign rom[13'h149e] = 0;
    assign rom[13'h149f] = 0;
    assign rom[13'h14a0] = 0;
    assign rom[13'h14a1] = 1;
    assign rom[13'h14a2] = 1;
    assign rom[13'h14a3] = 0;
    assign rom[13'h14a4] = 0;
    assign rom[13'h14a5] = 1;
    assign rom[13'h14a6] = 1;
    assign rom[13'h14a7] = 0;
    assign rom[13'h14a8] = 0;
    assign rom[13'h14a9] = 1;
    assign rom[13'h14aa] = 1;
    assign rom[13'h14ab] = 0;
    assign rom[13'h14ac] = 0;
    assign rom[13'h14ad] = 1;
    assign rom[13'h14ae] = 1;
    assign rom[13'h14af] = 0;
    assign rom[13'h14b0] = 0;
    assign rom[13'h14b1] = 1;
    assign rom[13'h14b2] = 1;
    assign rom[13'h14b3] = 0;
    assign rom[13'h14b4] = 0;
    assign rom[13'h14b5] = 1;
    assign rom[13'h14b6] = 1;
    assign rom[13'h14b7] = 0;
    assign rom[13'h14b8] = 0;
    assign rom[13'h14b9] = 0;
    assign rom[13'h14ba] = 0;
    assign rom[13'h14bb] = 0;
    assign rom[13'h14bc] = 0;
    assign rom[13'h14bd] = 0;
    assign rom[13'h14be] = 0;
    assign rom[13'h14bf] = 0;
    assign rom[13'h14c0] = 0;
    assign rom[13'h14c1] = 0;
    assign rom[13'h14c2] = 1;
    assign rom[13'h14c3] = 1;
    assign rom[13'h14c4] = 1;
    assign rom[13'h14c5] = 1;
    assign rom[13'h14c6] = 1;
    assign rom[13'h14c7] = 0;
    assign rom[13'h14c8] = 0;
    assign rom[13'h14c9] = 1;
    assign rom[13'h14ca] = 1;
    assign rom[13'h14cb] = 0;
    assign rom[13'h14cc] = 0;
    assign rom[13'h14cd] = 0;
    assign rom[13'h14ce] = 0;
    assign rom[13'h14cf] = 0;
    assign rom[13'h14d0] = 0;
    assign rom[13'h14d1] = 1;
    assign rom[13'h14d2] = 1;
    assign rom[13'h14d3] = 0;
    assign rom[13'h14d4] = 0;
    assign rom[13'h14d5] = 0;
    assign rom[13'h14d6] = 0;
    assign rom[13'h14d7] = 0;
    assign rom[13'h14d8] = 0;
    assign rom[13'h14d9] = 0;
    assign rom[13'h14da] = 1;
    assign rom[13'h14db] = 1;
    assign rom[13'h14dc] = 1;
    assign rom[13'h14dd] = 1;
    assign rom[13'h14de] = 0;
    assign rom[13'h14df] = 0;
    assign rom[13'h14e0] = 0;
    assign rom[13'h14e1] = 0;
    assign rom[13'h14e2] = 0;
    assign rom[13'h14e3] = 0;
    assign rom[13'h14e4] = 0;
    assign rom[13'h14e5] = 1;
    assign rom[13'h14e6] = 1;
    assign rom[13'h14e7] = 0;
    assign rom[13'h14e8] = 0;
    assign rom[13'h14e9] = 0;
    assign rom[13'h14ea] = 0;
    assign rom[13'h14eb] = 0;
    assign rom[13'h14ec] = 0;
    assign rom[13'h14ed] = 1;
    assign rom[13'h14ee] = 1;
    assign rom[13'h14ef] = 0;
    assign rom[13'h14f0] = 0;
    assign rom[13'h14f1] = 1;
    assign rom[13'h14f2] = 1;
    assign rom[13'h14f3] = 1;
    assign rom[13'h14f4] = 1;
    assign rom[13'h14f5] = 1;
    assign rom[13'h14f6] = 0;
    assign rom[13'h14f7] = 0;
    assign rom[13'h14f8] = 0;
    assign rom[13'h14f9] = 0;
    assign rom[13'h14fa] = 0;
    assign rom[13'h14fb] = 0;
    assign rom[13'h14fc] = 0;
    assign rom[13'h14fd] = 0;
    assign rom[13'h14fe] = 0;
    assign rom[13'h14ff] = 0;
    assign rom[13'h1500] = 0;
    assign rom[13'h1501] = 1;
    assign rom[13'h1502] = 1;
    assign rom[13'h1503] = 1;
    assign rom[13'h1504] = 1;
    assign rom[13'h1505] = 1;
    assign rom[13'h1506] = 1;
    assign rom[13'h1507] = 0;
    assign rom[13'h1508] = 0;
    assign rom[13'h1509] = 0;
    assign rom[13'h150a] = 0;
    assign rom[13'h150b] = 1;
    assign rom[13'h150c] = 1;
    assign rom[13'h150d] = 0;
    assign rom[13'h150e] = 0;
    assign rom[13'h150f] = 0;
    assign rom[13'h1510] = 0;
    assign rom[13'h1511] = 0;
    assign rom[13'h1512] = 0;
    assign rom[13'h1513] = 1;
    assign rom[13'h1514] = 1;
    assign rom[13'h1515] = 0;
    assign rom[13'h1516] = 0;
    assign rom[13'h1517] = 0;
    assign rom[13'h1518] = 0;
    assign rom[13'h1519] = 0;
    assign rom[13'h151a] = 0;
    assign rom[13'h151b] = 1;
    assign rom[13'h151c] = 1;
    assign rom[13'h151d] = 0;
    assign rom[13'h151e] = 0;
    assign rom[13'h151f] = 0;
    assign rom[13'h1520] = 0;
    assign rom[13'h1521] = 0;
    assign rom[13'h1522] = 0;
    assign rom[13'h1523] = 1;
    assign rom[13'h1524] = 1;
    assign rom[13'h1525] = 0;
    assign rom[13'h1526] = 0;
    assign rom[13'h1527] = 0;
    assign rom[13'h1528] = 0;
    assign rom[13'h1529] = 0;
    assign rom[13'h152a] = 0;
    assign rom[13'h152b] = 1;
    assign rom[13'h152c] = 1;
    assign rom[13'h152d] = 0;
    assign rom[13'h152e] = 0;
    assign rom[13'h152f] = 0;
    assign rom[13'h1530] = 0;
    assign rom[13'h1531] = 0;
    assign rom[13'h1532] = 0;
    assign rom[13'h1533] = 1;
    assign rom[13'h1534] = 1;
    assign rom[13'h1535] = 0;
    assign rom[13'h1536] = 0;
    assign rom[13'h1537] = 0;
    assign rom[13'h1538] = 0;
    assign rom[13'h1539] = 0;
    assign rom[13'h153a] = 0;
    assign rom[13'h153b] = 0;
    assign rom[13'h153c] = 0;
    assign rom[13'h153d] = 0;
    assign rom[13'h153e] = 0;
    assign rom[13'h153f] = 0;
    assign rom[13'h1540] = 0;
    assign rom[13'h1541] = 1;
    assign rom[13'h1542] = 1;
    assign rom[13'h1543] = 0;
    assign rom[13'h1544] = 0;
    assign rom[13'h1545] = 1;
    assign rom[13'h1546] = 1;
    assign rom[13'h1547] = 0;
    assign rom[13'h1548] = 0;
    assign rom[13'h1549] = 1;
    assign rom[13'h154a] = 1;
    assign rom[13'h154b] = 0;
    assign rom[13'h154c] = 0;
    assign rom[13'h154d] = 1;
    assign rom[13'h154e] = 1;
    assign rom[13'h154f] = 0;
    assign rom[13'h1550] = 0;
    assign rom[13'h1551] = 1;
    assign rom[13'h1552] = 1;
    assign rom[13'h1553] = 0;
    assign rom[13'h1554] = 0;
    assign rom[13'h1555] = 1;
    assign rom[13'h1556] = 1;
    assign rom[13'h1557] = 0;
    assign rom[13'h1558] = 0;
    assign rom[13'h1559] = 1;
    assign rom[13'h155a] = 1;
    assign rom[13'h155b] = 0;
    assign rom[13'h155c] = 0;
    assign rom[13'h155d] = 1;
    assign rom[13'h155e] = 1;
    assign rom[13'h155f] = 0;
    assign rom[13'h1560] = 0;
    assign rom[13'h1561] = 1;
    assign rom[13'h1562] = 1;
    assign rom[13'h1563] = 0;
    assign rom[13'h1564] = 0;
    assign rom[13'h1565] = 1;
    assign rom[13'h1566] = 1;
    assign rom[13'h1567] = 0;
    assign rom[13'h1568] = 0;
    assign rom[13'h1569] = 1;
    assign rom[13'h156a] = 1;
    assign rom[13'h156b] = 0;
    assign rom[13'h156c] = 0;
    assign rom[13'h156d] = 1;
    assign rom[13'h156e] = 1;
    assign rom[13'h156f] = 0;
    assign rom[13'h1570] = 0;
    assign rom[13'h1571] = 0;
    assign rom[13'h1572] = 1;
    assign rom[13'h1573] = 1;
    assign rom[13'h1574] = 1;
    assign rom[13'h1575] = 1;
    assign rom[13'h1576] = 0;
    assign rom[13'h1577] = 0;
    assign rom[13'h1578] = 0;
    assign rom[13'h1579] = 0;
    assign rom[13'h157a] = 0;
    assign rom[13'h157b] = 0;
    assign rom[13'h157c] = 0;
    assign rom[13'h157d] = 0;
    assign rom[13'h157e] = 0;
    assign rom[13'h157f] = 0;
    assign rom[13'h1580] = 0;
    assign rom[13'h1581] = 1;
    assign rom[13'h1582] = 1;
    assign rom[13'h1583] = 0;
    assign rom[13'h1584] = 0;
    assign rom[13'h1585] = 1;
    assign rom[13'h1586] = 1;
    assign rom[13'h1587] = 0;
    assign rom[13'h1588] = 0;
    assign rom[13'h1589] = 1;
    assign rom[13'h158a] = 1;
    assign rom[13'h158b] = 0;
    assign rom[13'h158c] = 0;
    assign rom[13'h158d] = 1;
    assign rom[13'h158e] = 1;
    assign rom[13'h158f] = 0;
    assign rom[13'h1590] = 0;
    assign rom[13'h1591] = 1;
    assign rom[13'h1592] = 1;
    assign rom[13'h1593] = 0;
    assign rom[13'h1594] = 0;
    assign rom[13'h1595] = 1;
    assign rom[13'h1596] = 1;
    assign rom[13'h1597] = 0;
    assign rom[13'h1598] = 0;
    assign rom[13'h1599] = 1;
    assign rom[13'h159a] = 1;
    assign rom[13'h159b] = 0;
    assign rom[13'h159c] = 0;
    assign rom[13'h159d] = 1;
    assign rom[13'h159e] = 1;
    assign rom[13'h159f] = 0;
    assign rom[13'h15a0] = 0;
    assign rom[13'h15a1] = 0;
    assign rom[13'h15a2] = 1;
    assign rom[13'h15a3] = 1;
    assign rom[13'h15a4] = 1;
    assign rom[13'h15a5] = 1;
    assign rom[13'h15a6] = 0;
    assign rom[13'h15a7] = 0;
    assign rom[13'h15a8] = 0;
    assign rom[13'h15a9] = 0;
    assign rom[13'h15aa] = 1;
    assign rom[13'h15ab] = 1;
    assign rom[13'h15ac] = 1;
    assign rom[13'h15ad] = 1;
    assign rom[13'h15ae] = 0;
    assign rom[13'h15af] = 0;
    assign rom[13'h15b0] = 0;
    assign rom[13'h15b1] = 0;
    assign rom[13'h15b2] = 0;
    assign rom[13'h15b3] = 1;
    assign rom[13'h15b4] = 1;
    assign rom[13'h15b5] = 0;
    assign rom[13'h15b6] = 0;
    assign rom[13'h15b7] = 0;
    assign rom[13'h15b8] = 0;
    assign rom[13'h15b9] = 0;
    assign rom[13'h15ba] = 0;
    assign rom[13'h15bb] = 0;
    assign rom[13'h15bc] = 0;
    assign rom[13'h15bd] = 0;
    assign rom[13'h15be] = 0;
    assign rom[13'h15bf] = 0;
    assign rom[13'h15c0] = 1;
    assign rom[13'h15c1] = 1;
    assign rom[13'h15c2] = 0;
    assign rom[13'h15c3] = 0;
    assign rom[13'h15c4] = 0;
    assign rom[13'h15c5] = 1;
    assign rom[13'h15c6] = 1;
    assign rom[13'h15c7] = 0;
    assign rom[13'h15c8] = 1;
    assign rom[13'h15c9] = 1;
    assign rom[13'h15ca] = 0;
    assign rom[13'h15cb] = 0;
    assign rom[13'h15cc] = 0;
    assign rom[13'h15cd] = 1;
    assign rom[13'h15ce] = 1;
    assign rom[13'h15cf] = 0;
    assign rom[13'h15d0] = 1;
    assign rom[13'h15d1] = 1;
    assign rom[13'h15d2] = 0;
    assign rom[13'h15d3] = 1;
    assign rom[13'h15d4] = 0;
    assign rom[13'h15d5] = 1;
    assign rom[13'h15d6] = 1;
    assign rom[13'h15d7] = 0;
    assign rom[13'h15d8] = 1;
    assign rom[13'h15d9] = 1;
    assign rom[13'h15da] = 0;
    assign rom[13'h15db] = 1;
    assign rom[13'h15dc] = 0;
    assign rom[13'h15dd] = 1;
    assign rom[13'h15de] = 1;
    assign rom[13'h15df] = 0;
    assign rom[13'h15e0] = 1;
    assign rom[13'h15e1] = 1;
    assign rom[13'h15e2] = 1;
    assign rom[13'h15e3] = 1;
    assign rom[13'h15e4] = 1;
    assign rom[13'h15e5] = 1;
    assign rom[13'h15e6] = 1;
    assign rom[13'h15e7] = 0;
    assign rom[13'h15e8] = 1;
    assign rom[13'h15e9] = 1;
    assign rom[13'h15ea] = 1;
    assign rom[13'h15eb] = 0;
    assign rom[13'h15ec] = 1;
    assign rom[13'h15ed] = 1;
    assign rom[13'h15ee] = 1;
    assign rom[13'h15ef] = 0;
    assign rom[13'h15f0] = 0;
    assign rom[13'h15f1] = 1;
    assign rom[13'h15f2] = 0;
    assign rom[13'h15f3] = 0;
    assign rom[13'h15f4] = 0;
    assign rom[13'h15f5] = 1;
    assign rom[13'h15f6] = 0;
    assign rom[13'h15f7] = 0;
    assign rom[13'h15f8] = 0;
    assign rom[13'h15f9] = 0;
    assign rom[13'h15fa] = 0;
    assign rom[13'h15fb] = 0;
    assign rom[13'h15fc] = 0;
    assign rom[13'h15fd] = 0;
    assign rom[13'h15fe] = 0;
    assign rom[13'h15ff] = 0;
    assign rom[13'h1600] = 0;
    assign rom[13'h1601] = 1;
    assign rom[13'h1602] = 1;
    assign rom[13'h1603] = 0;
    assign rom[13'h1604] = 0;
    assign rom[13'h1605] = 1;
    assign rom[13'h1606] = 1;
    assign rom[13'h1607] = 0;
    assign rom[13'h1608] = 0;
    assign rom[13'h1609] = 1;
    assign rom[13'h160a] = 1;
    assign rom[13'h160b] = 0;
    assign rom[13'h160c] = 0;
    assign rom[13'h160d] = 1;
    assign rom[13'h160e] = 1;
    assign rom[13'h160f] = 0;
    assign rom[13'h1610] = 0;
    assign rom[13'h1611] = 0;
    assign rom[13'h1612] = 1;
    assign rom[13'h1613] = 1;
    assign rom[13'h1614] = 1;
    assign rom[13'h1615] = 1;
    assign rom[13'h1616] = 0;
    assign rom[13'h1617] = 0;
    assign rom[13'h1618] = 0;
    assign rom[13'h1619] = 0;
    assign rom[13'h161a] = 0;
    assign rom[13'h161b] = 1;
    assign rom[13'h161c] = 1;
    assign rom[13'h161d] = 0;
    assign rom[13'h161e] = 0;
    assign rom[13'h161f] = 0;
    assign rom[13'h1620] = 0;
    assign rom[13'h1621] = 0;
    assign rom[13'h1622] = 1;
    assign rom[13'h1623] = 1;
    assign rom[13'h1624] = 1;
    assign rom[13'h1625] = 1;
    assign rom[13'h1626] = 0;
    assign rom[13'h1627] = 0;
    assign rom[13'h1628] = 0;
    assign rom[13'h1629] = 1;
    assign rom[13'h162a] = 1;
    assign rom[13'h162b] = 0;
    assign rom[13'h162c] = 0;
    assign rom[13'h162d] = 1;
    assign rom[13'h162e] = 1;
    assign rom[13'h162f] = 0;
    assign rom[13'h1630] = 0;
    assign rom[13'h1631] = 1;
    assign rom[13'h1632] = 1;
    assign rom[13'h1633] = 0;
    assign rom[13'h1634] = 0;
    assign rom[13'h1635] = 1;
    assign rom[13'h1636] = 1;
    assign rom[13'h1637] = 0;
    assign rom[13'h1638] = 0;
    assign rom[13'h1639] = 0;
    assign rom[13'h163a] = 0;
    assign rom[13'h163b] = 0;
    assign rom[13'h163c] = 0;
    assign rom[13'h163d] = 0;
    assign rom[13'h163e] = 0;
    assign rom[13'h163f] = 0;
    assign rom[13'h1640] = 0;
    assign rom[13'h1641] = 1;
    assign rom[13'h1642] = 1;
    assign rom[13'h1643] = 0;
    assign rom[13'h1644] = 0;
    assign rom[13'h1645] = 1;
    assign rom[13'h1646] = 1;
    assign rom[13'h1647] = 0;
    assign rom[13'h1648] = 0;
    assign rom[13'h1649] = 1;
    assign rom[13'h164a] = 1;
    assign rom[13'h164b] = 0;
    assign rom[13'h164c] = 0;
    assign rom[13'h164d] = 1;
    assign rom[13'h164e] = 1;
    assign rom[13'h164f] = 0;
    assign rom[13'h1650] = 0;
    assign rom[13'h1651] = 1;
    assign rom[13'h1652] = 1;
    assign rom[13'h1653] = 0;
    assign rom[13'h1654] = 0;
    assign rom[13'h1655] = 1;
    assign rom[13'h1656] = 1;
    assign rom[13'h1657] = 0;
    assign rom[13'h1658] = 0;
    assign rom[13'h1659] = 0;
    assign rom[13'h165a] = 1;
    assign rom[13'h165b] = 1;
    assign rom[13'h165c] = 1;
    assign rom[13'h165d] = 1;
    assign rom[13'h165e] = 0;
    assign rom[13'h165f] = 0;
    assign rom[13'h1660] = 0;
    assign rom[13'h1661] = 0;
    assign rom[13'h1662] = 0;
    assign rom[13'h1663] = 1;
    assign rom[13'h1664] = 1;
    assign rom[13'h1665] = 0;
    assign rom[13'h1666] = 0;
    assign rom[13'h1667] = 0;
    assign rom[13'h1668] = 0;
    assign rom[13'h1669] = 0;
    assign rom[13'h166a] = 0;
    assign rom[13'h166b] = 1;
    assign rom[13'h166c] = 1;
    assign rom[13'h166d] = 0;
    assign rom[13'h166e] = 0;
    assign rom[13'h166f] = 0;
    assign rom[13'h1670] = 0;
    assign rom[13'h1671] = 0;
    assign rom[13'h1672] = 0;
    assign rom[13'h1673] = 1;
    assign rom[13'h1674] = 1;
    assign rom[13'h1675] = 0;
    assign rom[13'h1676] = 0;
    assign rom[13'h1677] = 0;
    assign rom[13'h1678] = 0;
    assign rom[13'h1679] = 0;
    assign rom[13'h167a] = 0;
    assign rom[13'h167b] = 0;
    assign rom[13'h167c] = 0;
    assign rom[13'h167d] = 0;
    assign rom[13'h167e] = 0;
    assign rom[13'h167f] = 0;
    assign rom[13'h1680] = 0;
    assign rom[13'h1681] = 1;
    assign rom[13'h1682] = 1;
    assign rom[13'h1683] = 1;
    assign rom[13'h1684] = 1;
    assign rom[13'h1685] = 1;
    assign rom[13'h1686] = 1;
    assign rom[13'h1687] = 0;
    assign rom[13'h1688] = 0;
    assign rom[13'h1689] = 0;
    assign rom[13'h168a] = 0;
    assign rom[13'h168b] = 0;
    assign rom[13'h168c] = 0;
    assign rom[13'h168d] = 1;
    assign rom[13'h168e] = 1;
    assign rom[13'h168f] = 0;
    assign rom[13'h1690] = 0;
    assign rom[13'h1691] = 0;
    assign rom[13'h1692] = 0;
    assign rom[13'h1693] = 0;
    assign rom[13'h1694] = 1;
    assign rom[13'h1695] = 1;
    assign rom[13'h1696] = 0;
    assign rom[13'h1697] = 0;
    assign rom[13'h1698] = 0;
    assign rom[13'h1699] = 0;
    assign rom[13'h169a] = 0;
    assign rom[13'h169b] = 1;
    assign rom[13'h169c] = 1;
    assign rom[13'h169d] = 0;
    assign rom[13'h169e] = 0;
    assign rom[13'h169f] = 0;
    assign rom[13'h16a0] = 0;
    assign rom[13'h16a1] = 0;
    assign rom[13'h16a2] = 1;
    assign rom[13'h16a3] = 1;
    assign rom[13'h16a4] = 0;
    assign rom[13'h16a5] = 0;
    assign rom[13'h16a6] = 0;
    assign rom[13'h16a7] = 0;
    assign rom[13'h16a8] = 0;
    assign rom[13'h16a9] = 1;
    assign rom[13'h16aa] = 1;
    assign rom[13'h16ab] = 0;
    assign rom[13'h16ac] = 0;
    assign rom[13'h16ad] = 0;
    assign rom[13'h16ae] = 0;
    assign rom[13'h16af] = 0;
    assign rom[13'h16b0] = 0;
    assign rom[13'h16b1] = 1;
    assign rom[13'h16b2] = 1;
    assign rom[13'h16b3] = 1;
    assign rom[13'h16b4] = 1;
    assign rom[13'h16b5] = 1;
    assign rom[13'h16b6] = 1;
    assign rom[13'h16b7] = 0;
    assign rom[13'h16b8] = 0;
    assign rom[13'h16b9] = 0;
    assign rom[13'h16ba] = 0;
    assign rom[13'h16bb] = 0;
    assign rom[13'h16bc] = 0;
    assign rom[13'h16bd] = 0;
    assign rom[13'h16be] = 0;
    assign rom[13'h16bf] = 0;
    assign rom[13'h16c0] = 0;
    assign rom[13'h16c1] = 0;
    assign rom[13'h16c2] = 1;
    assign rom[13'h16c3] = 1;
    assign rom[13'h16c4] = 1;
    assign rom[13'h16c5] = 1;
    assign rom[13'h16c6] = 0;
    assign rom[13'h16c7] = 0;
    assign rom[13'h16c8] = 0;
    assign rom[13'h16c9] = 0;
    assign rom[13'h16ca] = 1;
    assign rom[13'h16cb] = 1;
    assign rom[13'h16cc] = 0;
    assign rom[13'h16cd] = 0;
    assign rom[13'h16ce] = 0;
    assign rom[13'h16cf] = 0;
    assign rom[13'h16d0] = 0;
    assign rom[13'h16d1] = 0;
    assign rom[13'h16d2] = 1;
    assign rom[13'h16d3] = 1;
    assign rom[13'h16d4] = 0;
    assign rom[13'h16d5] = 0;
    assign rom[13'h16d6] = 0;
    assign rom[13'h16d7] = 0;
    assign rom[13'h16d8] = 0;
    assign rom[13'h16d9] = 0;
    assign rom[13'h16da] = 1;
    assign rom[13'h16db] = 1;
    assign rom[13'h16dc] = 0;
    assign rom[13'h16dd] = 0;
    assign rom[13'h16de] = 0;
    assign rom[13'h16df] = 0;
    assign rom[13'h16e0] = 0;
    assign rom[13'h16e1] = 0;
    assign rom[13'h16e2] = 1;
    assign rom[13'h16e3] = 1;
    assign rom[13'h16e4] = 0;
    assign rom[13'h16e5] = 0;
    assign rom[13'h16e6] = 0;
    assign rom[13'h16e7] = 0;
    assign rom[13'h16e8] = 0;
    assign rom[13'h16e9] = 0;
    assign rom[13'h16ea] = 1;
    assign rom[13'h16eb] = 1;
    assign rom[13'h16ec] = 0;
    assign rom[13'h16ed] = 0;
    assign rom[13'h16ee] = 0;
    assign rom[13'h16ef] = 0;
    assign rom[13'h16f0] = 0;
    assign rom[13'h16f1] = 0;
    assign rom[13'h16f2] = 1;
    assign rom[13'h16f3] = 1;
    assign rom[13'h16f4] = 1;
    assign rom[13'h16f5] = 1;
    assign rom[13'h16f6] = 0;
    assign rom[13'h16f7] = 0;
    assign rom[13'h16f8] = 0;
    assign rom[13'h16f9] = 0;
    assign rom[13'h16fa] = 0;
    assign rom[13'h16fb] = 0;
    assign rom[13'h16fc] = 0;
    assign rom[13'h16fd] = 0;
    assign rom[13'h16fe] = 0;
    assign rom[13'h16ff] = 0;
    assign rom[13'h1700] = 0;
    assign rom[13'h1701] = 1;
    assign rom[13'h1702] = 0;
    assign rom[13'h1703] = 0;
    assign rom[13'h1704] = 0;
    assign rom[13'h1705] = 0;
    assign rom[13'h1706] = 0;
    assign rom[13'h1707] = 0;
    assign rom[13'h1708] = 0;
    assign rom[13'h1709] = 1;
    assign rom[13'h170a] = 1;
    assign rom[13'h170b] = 0;
    assign rom[13'h170c] = 0;
    assign rom[13'h170d] = 0;
    assign rom[13'h170e] = 0;
    assign rom[13'h170f] = 0;
    assign rom[13'h1710] = 0;
    assign rom[13'h1711] = 0;
    assign rom[13'h1712] = 1;
    assign rom[13'h1713] = 1;
    assign rom[13'h1714] = 0;
    assign rom[13'h1715] = 0;
    assign rom[13'h1716] = 0;
    assign rom[13'h1717] = 0;
    assign rom[13'h1718] = 0;
    assign rom[13'h1719] = 0;
    assign rom[13'h171a] = 0;
    assign rom[13'h171b] = 1;
    assign rom[13'h171c] = 1;
    assign rom[13'h171d] = 0;
    assign rom[13'h171e] = 0;
    assign rom[13'h171f] = 0;
    assign rom[13'h1720] = 0;
    assign rom[13'h1721] = 0;
    assign rom[13'h1722] = 0;
    assign rom[13'h1723] = 0;
    assign rom[13'h1724] = 1;
    assign rom[13'h1725] = 1;
    assign rom[13'h1726] = 0;
    assign rom[13'h1727] = 0;
    assign rom[13'h1728] = 0;
    assign rom[13'h1729] = 0;
    assign rom[13'h172a] = 0;
    assign rom[13'h172b] = 0;
    assign rom[13'h172c] = 0;
    assign rom[13'h172d] = 1;
    assign rom[13'h172e] = 1;
    assign rom[13'h172f] = 0;
    assign rom[13'h1730] = 0;
    assign rom[13'h1731] = 0;
    assign rom[13'h1732] = 0;
    assign rom[13'h1733] = 0;
    assign rom[13'h1734] = 0;
    assign rom[13'h1735] = 0;
    assign rom[13'h1736] = 1;
    assign rom[13'h1737] = 0;
    assign rom[13'h1738] = 0;
    assign rom[13'h1739] = 0;
    assign rom[13'h173a] = 0;
    assign rom[13'h173b] = 0;
    assign rom[13'h173c] = 0;
    assign rom[13'h173d] = 0;
    assign rom[13'h173e] = 0;
    assign rom[13'h173f] = 0;
    assign rom[13'h1740] = 0;
    assign rom[13'h1741] = 0;
    assign rom[13'h1742] = 1;
    assign rom[13'h1743] = 1;
    assign rom[13'h1744] = 1;
    assign rom[13'h1745] = 1;
    assign rom[13'h1746] = 0;
    assign rom[13'h1747] = 0;
    assign rom[13'h1748] = 0;
    assign rom[13'h1749] = 0;
    assign rom[13'h174a] = 0;
    assign rom[13'h174b] = 0;
    assign rom[13'h174c] = 1;
    assign rom[13'h174d] = 1;
    assign rom[13'h174e] = 0;
    assign rom[13'h174f] = 0;
    assign rom[13'h1750] = 0;
    assign rom[13'h1751] = 0;
    assign rom[13'h1752] = 0;
    assign rom[13'h1753] = 0;
    assign rom[13'h1754] = 1;
    assign rom[13'h1755] = 1;
    assign rom[13'h1756] = 0;
    assign rom[13'h1757] = 0;
    assign rom[13'h1758] = 0;
    assign rom[13'h1759] = 0;
    assign rom[13'h175a] = 0;
    assign rom[13'h175b] = 0;
    assign rom[13'h175c] = 1;
    assign rom[13'h175d] = 1;
    assign rom[13'h175e] = 0;
    assign rom[13'h175f] = 0;
    assign rom[13'h1760] = 0;
    assign rom[13'h1761] = 0;
    assign rom[13'h1762] = 0;
    assign rom[13'h1763] = 0;
    assign rom[13'h1764] = 1;
    assign rom[13'h1765] = 1;
    assign rom[13'h1766] = 0;
    assign rom[13'h1767] = 0;
    assign rom[13'h1768] = 0;
    assign rom[13'h1769] = 0;
    assign rom[13'h176a] = 0;
    assign rom[13'h176b] = 0;
    assign rom[13'h176c] = 1;
    assign rom[13'h176d] = 1;
    assign rom[13'h176e] = 0;
    assign rom[13'h176f] = 0;
    assign rom[13'h1770] = 0;
    assign rom[13'h1771] = 0;
    assign rom[13'h1772] = 1;
    assign rom[13'h1773] = 1;
    assign rom[13'h1774] = 1;
    assign rom[13'h1775] = 1;
    assign rom[13'h1776] = 0;
    assign rom[13'h1777] = 0;
    assign rom[13'h1778] = 0;
    assign rom[13'h1779] = 0;
    assign rom[13'h177a] = 0;
    assign rom[13'h177b] = 0;
    assign rom[13'h177c] = 0;
    assign rom[13'h177d] = 0;
    assign rom[13'h177e] = 0;
    assign rom[13'h177f] = 0;
    assign rom[13'h1780] = 0;
    assign rom[13'h1781] = 0;
    assign rom[13'h1782] = 0;
    assign rom[13'h1783] = 1;
    assign rom[13'h1784] = 0;
    assign rom[13'h1785] = 0;
    assign rom[13'h1786] = 0;
    assign rom[13'h1787] = 0;
    assign rom[13'h1788] = 0;
    assign rom[13'h1789] = 0;
    assign rom[13'h178a] = 1;
    assign rom[13'h178b] = 1;
    assign rom[13'h178c] = 1;
    assign rom[13'h178d] = 0;
    assign rom[13'h178e] = 0;
    assign rom[13'h178f] = 0;
    assign rom[13'h1790] = 0;
    assign rom[13'h1791] = 1;
    assign rom[13'h1792] = 1;
    assign rom[13'h1793] = 0;
    assign rom[13'h1794] = 1;
    assign rom[13'h1795] = 1;
    assign rom[13'h1796] = 0;
    assign rom[13'h1797] = 0;
    assign rom[13'h1798] = 0;
    assign rom[13'h1799] = 0;
    assign rom[13'h179a] = 0;
    assign rom[13'h179b] = 0;
    assign rom[13'h179c] = 0;
    assign rom[13'h179d] = 0;
    assign rom[13'h179e] = 0;
    assign rom[13'h179f] = 0;
    assign rom[13'h17a0] = 0;
    assign rom[13'h17a1] = 0;
    assign rom[13'h17a2] = 0;
    assign rom[13'h17a3] = 0;
    assign rom[13'h17a4] = 0;
    assign rom[13'h17a5] = 0;
    assign rom[13'h17a6] = 0;
    assign rom[13'h17a7] = 0;
    assign rom[13'h17a8] = 0;
    assign rom[13'h17a9] = 0;
    assign rom[13'h17aa] = 0;
    assign rom[13'h17ab] = 0;
    assign rom[13'h17ac] = 0;
    assign rom[13'h17ad] = 0;
    assign rom[13'h17ae] = 0;
    assign rom[13'h17af] = 0;
    assign rom[13'h17b0] = 0;
    assign rom[13'h17b1] = 0;
    assign rom[13'h17b2] = 0;
    assign rom[13'h17b3] = 0;
    assign rom[13'h17b4] = 0;
    assign rom[13'h17b5] = 0;
    assign rom[13'h17b6] = 0;
    assign rom[13'h17b7] = 0;
    assign rom[13'h17b8] = 0;
    assign rom[13'h17b9] = 0;
    assign rom[13'h17ba] = 0;
    assign rom[13'h17bb] = 0;
    assign rom[13'h17bc] = 0;
    assign rom[13'h17bd] = 0;
    assign rom[13'h17be] = 0;
    assign rom[13'h17bf] = 0;
    assign rom[13'h17c0] = 0;
    assign rom[13'h17c1] = 0;
    assign rom[13'h17c2] = 0;
    assign rom[13'h17c3] = 0;
    assign rom[13'h17c4] = 0;
    assign rom[13'h17c5] = 0;
    assign rom[13'h17c6] = 0;
    assign rom[13'h17c7] = 0;
    assign rom[13'h17c8] = 0;
    assign rom[13'h17c9] = 0;
    assign rom[13'h17ca] = 0;
    assign rom[13'h17cb] = 0;
    assign rom[13'h17cc] = 0;
    assign rom[13'h17cd] = 0;
    assign rom[13'h17ce] = 0;
    assign rom[13'h17cf] = 0;
    assign rom[13'h17d0] = 0;
    assign rom[13'h17d1] = 0;
    assign rom[13'h17d2] = 0;
    assign rom[13'h17d3] = 0;
    assign rom[13'h17d4] = 0;
    assign rom[13'h17d5] = 0;
    assign rom[13'h17d6] = 0;
    assign rom[13'h17d7] = 0;
    assign rom[13'h17d8] = 0;
    assign rom[13'h17d9] = 0;
    assign rom[13'h17da] = 0;
    assign rom[13'h17db] = 0;
    assign rom[13'h17dc] = 0;
    assign rom[13'h17dd] = 0;
    assign rom[13'h17de] = 0;
    assign rom[13'h17df] = 0;
    assign rom[13'h17e0] = 0;
    assign rom[13'h17e1] = 0;
    assign rom[13'h17e2] = 0;
    assign rom[13'h17e3] = 0;
    assign rom[13'h17e4] = 0;
    assign rom[13'h17e5] = 0;
    assign rom[13'h17e6] = 0;
    assign rom[13'h17e7] = 0;
    assign rom[13'h17e8] = 0;
    assign rom[13'h17e9] = 0;
    assign rom[13'h17ea] = 0;
    assign rom[13'h17eb] = 0;
    assign rom[13'h17ec] = 0;
    assign rom[13'h17ed] = 0;
    assign rom[13'h17ee] = 0;
    assign rom[13'h17ef] = 0;
    assign rom[13'h17f0] = 0;
    assign rom[13'h17f1] = 0;
    assign rom[13'h17f2] = 0;
    assign rom[13'h17f3] = 0;
    assign rom[13'h17f4] = 0;
    assign rom[13'h17f5] = 0;
    assign rom[13'h17f6] = 0;
    assign rom[13'h17f7] = 0;
    assign rom[13'h17f8] = 1;
    assign rom[13'h17f9] = 1;
    assign rom[13'h17fa] = 1;
    assign rom[13'h17fb] = 1;
    assign rom[13'h17fc] = 1;
    assign rom[13'h17fd] = 1;
    assign rom[13'h17fe] = 1;
    assign rom[13'h17ff] = 1;
    assign rom[13'h1800] = 0;
    assign rom[13'h1801] = 0;
    assign rom[13'h1802] = 0;
    assign rom[13'h1803] = 1;
    assign rom[13'h1804] = 1;
    assign rom[13'h1805] = 0;
    assign rom[13'h1806] = 0;
    assign rom[13'h1807] = 0;
    assign rom[13'h1808] = 0;
    assign rom[13'h1809] = 0;
    assign rom[13'h180a] = 0;
    assign rom[13'h180b] = 1;
    assign rom[13'h180c] = 1;
    assign rom[13'h180d] = 0;
    assign rom[13'h180e] = 0;
    assign rom[13'h180f] = 0;
    assign rom[13'h1810] = 0;
    assign rom[13'h1811] = 0;
    assign rom[13'h1812] = 0;
    assign rom[13'h1813] = 0;
    assign rom[13'h1814] = 1;
    assign rom[13'h1815] = 1;
    assign rom[13'h1816] = 0;
    assign rom[13'h1817] = 0;
    assign rom[13'h1818] = 0;
    assign rom[13'h1819] = 0;
    assign rom[13'h181a] = 0;
    assign rom[13'h181b] = 0;
    assign rom[13'h181c] = 0;
    assign rom[13'h181d] = 0;
    assign rom[13'h181e] = 0;
    assign rom[13'h181f] = 0;
    assign rom[13'h1820] = 0;
    assign rom[13'h1821] = 0;
    assign rom[13'h1822] = 0;
    assign rom[13'h1823] = 0;
    assign rom[13'h1824] = 0;
    assign rom[13'h1825] = 0;
    assign rom[13'h1826] = 0;
    assign rom[13'h1827] = 0;
    assign rom[13'h1828] = 0;
    assign rom[13'h1829] = 0;
    assign rom[13'h182a] = 0;
    assign rom[13'h182b] = 0;
    assign rom[13'h182c] = 0;
    assign rom[13'h182d] = 0;
    assign rom[13'h182e] = 0;
    assign rom[13'h182f] = 0;
    assign rom[13'h1830] = 0;
    assign rom[13'h1831] = 0;
    assign rom[13'h1832] = 0;
    assign rom[13'h1833] = 0;
    assign rom[13'h1834] = 0;
    assign rom[13'h1835] = 0;
    assign rom[13'h1836] = 0;
    assign rom[13'h1837] = 0;
    assign rom[13'h1838] = 0;
    assign rom[13'h1839] = 0;
    assign rom[13'h183a] = 0;
    assign rom[13'h183b] = 0;
    assign rom[13'h183c] = 0;
    assign rom[13'h183d] = 0;
    assign rom[13'h183e] = 0;
    assign rom[13'h183f] = 0;
    assign rom[13'h1840] = 0;
    assign rom[13'h1841] = 0;
    assign rom[13'h1842] = 0;
    assign rom[13'h1843] = 0;
    assign rom[13'h1844] = 0;
    assign rom[13'h1845] = 0;
    assign rom[13'h1846] = 0;
    assign rom[13'h1847] = 0;
    assign rom[13'h1848] = 0;
    assign rom[13'h1849] = 0;
    assign rom[13'h184a] = 0;
    assign rom[13'h184b] = 0;
    assign rom[13'h184c] = 0;
    assign rom[13'h184d] = 0;
    assign rom[13'h184e] = 0;
    assign rom[13'h184f] = 0;
    assign rom[13'h1850] = 0;
    assign rom[13'h1851] = 0;
    assign rom[13'h1852] = 1;
    assign rom[13'h1853] = 1;
    assign rom[13'h1854] = 1;
    assign rom[13'h1855] = 1;
    assign rom[13'h1856] = 0;
    assign rom[13'h1857] = 0;
    assign rom[13'h1858] = 0;
    assign rom[13'h1859] = 0;
    assign rom[13'h185a] = 0;
    assign rom[13'h185b] = 0;
    assign rom[13'h185c] = 0;
    assign rom[13'h185d] = 1;
    assign rom[13'h185e] = 1;
    assign rom[13'h185f] = 0;
    assign rom[13'h1860] = 0;
    assign rom[13'h1861] = 0;
    assign rom[13'h1862] = 1;
    assign rom[13'h1863] = 1;
    assign rom[13'h1864] = 1;
    assign rom[13'h1865] = 1;
    assign rom[13'h1866] = 1;
    assign rom[13'h1867] = 0;
    assign rom[13'h1868] = 0;
    assign rom[13'h1869] = 1;
    assign rom[13'h186a] = 1;
    assign rom[13'h186b] = 0;
    assign rom[13'h186c] = 0;
    assign rom[13'h186d] = 1;
    assign rom[13'h186e] = 1;
    assign rom[13'h186f] = 0;
    assign rom[13'h1870] = 0;
    assign rom[13'h1871] = 0;
    assign rom[13'h1872] = 1;
    assign rom[13'h1873] = 1;
    assign rom[13'h1874] = 1;
    assign rom[13'h1875] = 0;
    assign rom[13'h1876] = 1;
    assign rom[13'h1877] = 0;
    assign rom[13'h1878] = 0;
    assign rom[13'h1879] = 0;
    assign rom[13'h187a] = 0;
    assign rom[13'h187b] = 0;
    assign rom[13'h187c] = 0;
    assign rom[13'h187d] = 0;
    assign rom[13'h187e] = 0;
    assign rom[13'h187f] = 0;
    assign rom[13'h1880] = 0;
    assign rom[13'h1881] = 1;
    assign rom[13'h1882] = 1;
    assign rom[13'h1883] = 0;
    assign rom[13'h1884] = 0;
    assign rom[13'h1885] = 0;
    assign rom[13'h1886] = 0;
    assign rom[13'h1887] = 0;
    assign rom[13'h1888] = 0;
    assign rom[13'h1889] = 1;
    assign rom[13'h188a] = 1;
    assign rom[13'h188b] = 0;
    assign rom[13'h188c] = 0;
    assign rom[13'h188d] = 0;
    assign rom[13'h188e] = 0;
    assign rom[13'h188f] = 0;
    assign rom[13'h1890] = 0;
    assign rom[13'h1891] = 1;
    assign rom[13'h1892] = 1;
    assign rom[13'h1893] = 1;
    assign rom[13'h1894] = 1;
    assign rom[13'h1895] = 1;
    assign rom[13'h1896] = 0;
    assign rom[13'h1897] = 0;
    assign rom[13'h1898] = 0;
    assign rom[13'h1899] = 1;
    assign rom[13'h189a] = 1;
    assign rom[13'h189b] = 0;
    assign rom[13'h189c] = 0;
    assign rom[13'h189d] = 1;
    assign rom[13'h189e] = 1;
    assign rom[13'h189f] = 0;
    assign rom[13'h18a0] = 0;
    assign rom[13'h18a1] = 1;
    assign rom[13'h18a2] = 1;
    assign rom[13'h18a3] = 0;
    assign rom[13'h18a4] = 0;
    assign rom[13'h18a5] = 1;
    assign rom[13'h18a6] = 1;
    assign rom[13'h18a7] = 0;
    assign rom[13'h18a8] = 0;
    assign rom[13'h18a9] = 1;
    assign rom[13'h18aa] = 1;
    assign rom[13'h18ab] = 0;
    assign rom[13'h18ac] = 0;
    assign rom[13'h18ad] = 1;
    assign rom[13'h18ae] = 1;
    assign rom[13'h18af] = 0;
    assign rom[13'h18b0] = 0;
    assign rom[13'h18b1] = 1;
    assign rom[13'h18b2] = 1;
    assign rom[13'h18b3] = 1;
    assign rom[13'h18b4] = 1;
    assign rom[13'h18b5] = 1;
    assign rom[13'h18b6] = 0;
    assign rom[13'h18b7] = 0;
    assign rom[13'h18b8] = 0;
    assign rom[13'h18b9] = 0;
    assign rom[13'h18ba] = 0;
    assign rom[13'h18bb] = 0;
    assign rom[13'h18bc] = 0;
    assign rom[13'h18bd] = 0;
    assign rom[13'h18be] = 0;
    assign rom[13'h18bf] = 0;
    assign rom[13'h18c0] = 0;
    assign rom[13'h18c1] = 0;
    assign rom[13'h18c2] = 0;
    assign rom[13'h18c3] = 0;
    assign rom[13'h18c4] = 0;
    assign rom[13'h18c5] = 0;
    assign rom[13'h18c6] = 0;
    assign rom[13'h18c7] = 0;
    assign rom[13'h18c8] = 0;
    assign rom[13'h18c9] = 0;
    assign rom[13'h18ca] = 0;
    assign rom[13'h18cb] = 0;
    assign rom[13'h18cc] = 0;
    assign rom[13'h18cd] = 0;
    assign rom[13'h18ce] = 0;
    assign rom[13'h18cf] = 0;
    assign rom[13'h18d0] = 0;
    assign rom[13'h18d1] = 0;
    assign rom[13'h18d2] = 1;
    assign rom[13'h18d3] = 1;
    assign rom[13'h18d4] = 1;
    assign rom[13'h18d5] = 1;
    assign rom[13'h18d6] = 0;
    assign rom[13'h18d7] = 0;
    assign rom[13'h18d8] = 0;
    assign rom[13'h18d9] = 1;
    assign rom[13'h18da] = 1;
    assign rom[13'h18db] = 0;
    assign rom[13'h18dc] = 0;
    assign rom[13'h18dd] = 1;
    assign rom[13'h18de] = 1;
    assign rom[13'h18df] = 0;
    assign rom[13'h18e0] = 0;
    assign rom[13'h18e1] = 1;
    assign rom[13'h18e2] = 1;
    assign rom[13'h18e3] = 0;
    assign rom[13'h18e4] = 0;
    assign rom[13'h18e5] = 0;
    assign rom[13'h18e6] = 0;
    assign rom[13'h18e7] = 0;
    assign rom[13'h18e8] = 0;
    assign rom[13'h18e9] = 1;
    assign rom[13'h18ea] = 1;
    assign rom[13'h18eb] = 0;
    assign rom[13'h18ec] = 0;
    assign rom[13'h18ed] = 1;
    assign rom[13'h18ee] = 1;
    assign rom[13'h18ef] = 0;
    assign rom[13'h18f0] = 0;
    assign rom[13'h18f1] = 0;
    assign rom[13'h18f2] = 1;
    assign rom[13'h18f3] = 1;
    assign rom[13'h18f4] = 1;
    assign rom[13'h18f5] = 1;
    assign rom[13'h18f6] = 0;
    assign rom[13'h18f7] = 0;
    assign rom[13'h18f8] = 0;
    assign rom[13'h18f9] = 0;
    assign rom[13'h18fa] = 0;
    assign rom[13'h18fb] = 0;
    assign rom[13'h18fc] = 0;
    assign rom[13'h18fd] = 0;
    assign rom[13'h18fe] = 0;
    assign rom[13'h18ff] = 0;
    assign rom[13'h1900] = 0;
    assign rom[13'h1901] = 0;
    assign rom[13'h1902] = 0;
    assign rom[13'h1903] = 0;
    assign rom[13'h1904] = 0;
    assign rom[13'h1905] = 1;
    assign rom[13'h1906] = 1;
    assign rom[13'h1907] = 0;
    assign rom[13'h1908] = 0;
    assign rom[13'h1909] = 0;
    assign rom[13'h190a] = 0;
    assign rom[13'h190b] = 0;
    assign rom[13'h190c] = 0;
    assign rom[13'h190d] = 1;
    assign rom[13'h190e] = 1;
    assign rom[13'h190f] = 0;
    assign rom[13'h1910] = 0;
    assign rom[13'h1911] = 0;
    assign rom[13'h1912] = 1;
    assign rom[13'h1913] = 1;
    assign rom[13'h1914] = 1;
    assign rom[13'h1915] = 1;
    assign rom[13'h1916] = 1;
    assign rom[13'h1917] = 0;
    assign rom[13'h1918] = 0;
    assign rom[13'h1919] = 1;
    assign rom[13'h191a] = 1;
    assign rom[13'h191b] = 0;
    assign rom[13'h191c] = 0;
    assign rom[13'h191d] = 1;
    assign rom[13'h191e] = 1;
    assign rom[13'h191f] = 0;
    assign rom[13'h1920] = 0;
    assign rom[13'h1921] = 1;
    assign rom[13'h1922] = 1;
    assign rom[13'h1923] = 0;
    assign rom[13'h1924] = 0;
    assign rom[13'h1925] = 1;
    assign rom[13'h1926] = 1;
    assign rom[13'h1927] = 0;
    assign rom[13'h1928] = 0;
    assign rom[13'h1929] = 1;
    assign rom[13'h192a] = 1;
    assign rom[13'h192b] = 0;
    assign rom[13'h192c] = 0;
    assign rom[13'h192d] = 1;
    assign rom[13'h192e] = 1;
    assign rom[13'h192f] = 0;
    assign rom[13'h1930] = 0;
    assign rom[13'h1931] = 0;
    assign rom[13'h1932] = 1;
    assign rom[13'h1933] = 1;
    assign rom[13'h1934] = 1;
    assign rom[13'h1935] = 1;
    assign rom[13'h1936] = 1;
    assign rom[13'h1937] = 0;
    assign rom[13'h1938] = 0;
    assign rom[13'h1939] = 0;
    assign rom[13'h193a] = 0;
    assign rom[13'h193b] = 0;
    assign rom[13'h193c] = 0;
    assign rom[13'h193d] = 0;
    assign rom[13'h193e] = 0;
    assign rom[13'h193f] = 0;
    assign rom[13'h1940] = 0;
    assign rom[13'h1941] = 0;
    assign rom[13'h1942] = 0;
    assign rom[13'h1943] = 0;
    assign rom[13'h1944] = 0;
    assign rom[13'h1945] = 0;
    assign rom[13'h1946] = 0;
    assign rom[13'h1947] = 0;
    assign rom[13'h1948] = 0;
    assign rom[13'h1949] = 0;
    assign rom[13'h194a] = 0;
    assign rom[13'h194b] = 0;
    assign rom[13'h194c] = 0;
    assign rom[13'h194d] = 0;
    assign rom[13'h194e] = 0;
    assign rom[13'h194f] = 0;
    assign rom[13'h1950] = 0;
    assign rom[13'h1951] = 0;
    assign rom[13'h1952] = 1;
    assign rom[13'h1953] = 1;
    assign rom[13'h1954] = 1;
    assign rom[13'h1955] = 1;
    assign rom[13'h1956] = 0;
    assign rom[13'h1957] = 0;
    assign rom[13'h1958] = 0;
    assign rom[13'h1959] = 1;
    assign rom[13'h195a] = 1;
    assign rom[13'h195b] = 0;
    assign rom[13'h195c] = 0;
    assign rom[13'h195d] = 1;
    assign rom[13'h195e] = 1;
    assign rom[13'h195f] = 0;
    assign rom[13'h1960] = 0;
    assign rom[13'h1961] = 1;
    assign rom[13'h1962] = 1;
    assign rom[13'h1963] = 1;
    assign rom[13'h1964] = 1;
    assign rom[13'h1965] = 1;
    assign rom[13'h1966] = 0;
    assign rom[13'h1967] = 0;
    assign rom[13'h1968] = 0;
    assign rom[13'h1969] = 1;
    assign rom[13'h196a] = 1;
    assign rom[13'h196b] = 0;
    assign rom[13'h196c] = 0;
    assign rom[13'h196d] = 0;
    assign rom[13'h196e] = 0;
    assign rom[13'h196f] = 0;
    assign rom[13'h1970] = 0;
    assign rom[13'h1971] = 0;
    assign rom[13'h1972] = 1;
    assign rom[13'h1973] = 1;
    assign rom[13'h1974] = 1;
    assign rom[13'h1975] = 1;
    assign rom[13'h1976] = 0;
    assign rom[13'h1977] = 0;
    assign rom[13'h1978] = 0;
    assign rom[13'h1979] = 0;
    assign rom[13'h197a] = 0;
    assign rom[13'h197b] = 0;
    assign rom[13'h197c] = 0;
    assign rom[13'h197d] = 0;
    assign rom[13'h197e] = 0;
    assign rom[13'h197f] = 0;
    assign rom[13'h1980] = 0;
    assign rom[13'h1981] = 0;
    assign rom[13'h1982] = 0;
    assign rom[13'h1983] = 0;
    assign rom[13'h1984] = 1;
    assign rom[13'h1985] = 1;
    assign rom[13'h1986] = 1;
    assign rom[13'h1987] = 0;
    assign rom[13'h1988] = 0;
    assign rom[13'h1989] = 0;
    assign rom[13'h198a] = 0;
    assign rom[13'h198b] = 1;
    assign rom[13'h198c] = 1;
    assign rom[13'h198d] = 0;
    assign rom[13'h198e] = 0;
    assign rom[13'h198f] = 0;
    assign rom[13'h1990] = 0;
    assign rom[13'h1991] = 0;
    assign rom[13'h1992] = 0;
    assign rom[13'h1993] = 1;
    assign rom[13'h1994] = 1;
    assign rom[13'h1995] = 0;
    assign rom[13'h1996] = 0;
    assign rom[13'h1997] = 0;
    assign rom[13'h1998] = 0;
    assign rom[13'h1999] = 0;
    assign rom[13'h199a] = 1;
    assign rom[13'h199b] = 1;
    assign rom[13'h199c] = 1;
    assign rom[13'h199d] = 1;
    assign rom[13'h199e] = 1;
    assign rom[13'h199f] = 0;
    assign rom[13'h19a0] = 0;
    assign rom[13'h19a1] = 0;
    assign rom[13'h19a2] = 0;
    assign rom[13'h19a3] = 1;
    assign rom[13'h19a4] = 1;
    assign rom[13'h19a5] = 0;
    assign rom[13'h19a6] = 0;
    assign rom[13'h19a7] = 0;
    assign rom[13'h19a8] = 0;
    assign rom[13'h19a9] = 0;
    assign rom[13'h19aa] = 0;
    assign rom[13'h19ab] = 1;
    assign rom[13'h19ac] = 1;
    assign rom[13'h19ad] = 0;
    assign rom[13'h19ae] = 0;
    assign rom[13'h19af] = 0;
    assign rom[13'h19b0] = 0;
    assign rom[13'h19b1] = 0;
    assign rom[13'h19b2] = 0;
    assign rom[13'h19b3] = 1;
    assign rom[13'h19b4] = 1;
    assign rom[13'h19b5] = 0;
    assign rom[13'h19b6] = 0;
    assign rom[13'h19b7] = 0;
    assign rom[13'h19b8] = 0;
    assign rom[13'h19b9] = 0;
    assign rom[13'h19ba] = 0;
    assign rom[13'h19bb] = 0;
    assign rom[13'h19bc] = 0;
    assign rom[13'h19bd] = 0;
    assign rom[13'h19be] = 0;
    assign rom[13'h19bf] = 0;
    assign rom[13'h19c0] = 0;
    assign rom[13'h19c1] = 0;
    assign rom[13'h19c2] = 0;
    assign rom[13'h19c3] = 0;
    assign rom[13'h19c4] = 0;
    assign rom[13'h19c5] = 0;
    assign rom[13'h19c6] = 0;
    assign rom[13'h19c7] = 0;
    assign rom[13'h19c8] = 0;
    assign rom[13'h19c9] = 0;
    assign rom[13'h19ca] = 0;
    assign rom[13'h19cb] = 0;
    assign rom[13'h19cc] = 0;
    assign rom[13'h19cd] = 0;
    assign rom[13'h19ce] = 0;
    assign rom[13'h19cf] = 0;
    assign rom[13'h19d0] = 0;
    assign rom[13'h19d1] = 0;
    assign rom[13'h19d2] = 1;
    assign rom[13'h19d3] = 1;
    assign rom[13'h19d4] = 1;
    assign rom[13'h19d5] = 1;
    assign rom[13'h19d6] = 1;
    assign rom[13'h19d7] = 0;
    assign rom[13'h19d8] = 0;
    assign rom[13'h19d9] = 1;
    assign rom[13'h19da] = 1;
    assign rom[13'h19db] = 0;
    assign rom[13'h19dc] = 0;
    assign rom[13'h19dd] = 1;
    assign rom[13'h19de] = 1;
    assign rom[13'h19df] = 0;
    assign rom[13'h19e0] = 0;
    assign rom[13'h19e1] = 1;
    assign rom[13'h19e2] = 1;
    assign rom[13'h19e3] = 0;
    assign rom[13'h19e4] = 0;
    assign rom[13'h19e5] = 1;
    assign rom[13'h19e6] = 1;
    assign rom[13'h19e7] = 0;
    assign rom[13'h19e8] = 0;
    assign rom[13'h19e9] = 0;
    assign rom[13'h19ea] = 1;
    assign rom[13'h19eb] = 1;
    assign rom[13'h19ec] = 1;
    assign rom[13'h19ed] = 1;
    assign rom[13'h19ee] = 1;
    assign rom[13'h19ef] = 0;
    assign rom[13'h19f0] = 0;
    assign rom[13'h19f1] = 0;
    assign rom[13'h19f2] = 0;
    assign rom[13'h19f3] = 0;
    assign rom[13'h19f4] = 0;
    assign rom[13'h19f5] = 1;
    assign rom[13'h19f6] = 1;
    assign rom[13'h19f7] = 0;
    assign rom[13'h19f8] = 0;
    assign rom[13'h19f9] = 0;
    assign rom[13'h19fa] = 1;
    assign rom[13'h19fb] = 1;
    assign rom[13'h19fc] = 1;
    assign rom[13'h19fd] = 1;
    assign rom[13'h19fe] = 0;
    assign rom[13'h19ff] = 0;
    assign rom[13'h1a00] = 0;
    assign rom[13'h1a01] = 1;
    assign rom[13'h1a02] = 1;
    assign rom[13'h1a03] = 0;
    assign rom[13'h1a04] = 0;
    assign rom[13'h1a05] = 0;
    assign rom[13'h1a06] = 0;
    assign rom[13'h1a07] = 0;
    assign rom[13'h1a08] = 0;
    assign rom[13'h1a09] = 1;
    assign rom[13'h1a0a] = 1;
    assign rom[13'h1a0b] = 0;
    assign rom[13'h1a0c] = 0;
    assign rom[13'h1a0d] = 0;
    assign rom[13'h1a0e] = 0;
    assign rom[13'h1a0f] = 0;
    assign rom[13'h1a10] = 0;
    assign rom[13'h1a11] = 1;
    assign rom[13'h1a12] = 1;
    assign rom[13'h1a13] = 1;
    assign rom[13'h1a14] = 1;
    assign rom[13'h1a15] = 1;
    assign rom[13'h1a16] = 0;
    assign rom[13'h1a17] = 0;
    assign rom[13'h1a18] = 0;
    assign rom[13'h1a19] = 1;
    assign rom[13'h1a1a] = 1;
    assign rom[13'h1a1b] = 0;
    assign rom[13'h1a1c] = 0;
    assign rom[13'h1a1d] = 1;
    assign rom[13'h1a1e] = 1;
    assign rom[13'h1a1f] = 0;
    assign rom[13'h1a20] = 0;
    assign rom[13'h1a21] = 1;
    assign rom[13'h1a22] = 1;
    assign rom[13'h1a23] = 0;
    assign rom[13'h1a24] = 0;
    assign rom[13'h1a25] = 1;
    assign rom[13'h1a26] = 1;
    assign rom[13'h1a27] = 0;
    assign rom[13'h1a28] = 0;
    assign rom[13'h1a29] = 1;
    assign rom[13'h1a2a] = 1;
    assign rom[13'h1a2b] = 0;
    assign rom[13'h1a2c] = 0;
    assign rom[13'h1a2d] = 1;
    assign rom[13'h1a2e] = 1;
    assign rom[13'h1a2f] = 0;
    assign rom[13'h1a30] = 0;
    assign rom[13'h1a31] = 1;
    assign rom[13'h1a32] = 1;
    assign rom[13'h1a33] = 0;
    assign rom[13'h1a34] = 0;
    assign rom[13'h1a35] = 1;
    assign rom[13'h1a36] = 1;
    assign rom[13'h1a37] = 0;
    assign rom[13'h1a38] = 0;
    assign rom[13'h1a39] = 0;
    assign rom[13'h1a3a] = 0;
    assign rom[13'h1a3b] = 0;
    assign rom[13'h1a3c] = 0;
    assign rom[13'h1a3d] = 0;
    assign rom[13'h1a3e] = 0;
    assign rom[13'h1a3f] = 0;
    assign rom[13'h1a40] = 0;
    assign rom[13'h1a41] = 0;
    assign rom[13'h1a42] = 0;
    assign rom[13'h1a43] = 1;
    assign rom[13'h1a44] = 1;
    assign rom[13'h1a45] = 0;
    assign rom[13'h1a46] = 0;
    assign rom[13'h1a47] = 0;
    assign rom[13'h1a48] = 0;
    assign rom[13'h1a49] = 0;
    assign rom[13'h1a4a] = 0;
    assign rom[13'h1a4b] = 0;
    assign rom[13'h1a4c] = 0;
    assign rom[13'h1a4d] = 0;
    assign rom[13'h1a4e] = 0;
    assign rom[13'h1a4f] = 0;
    assign rom[13'h1a50] = 0;
    assign rom[13'h1a51] = 0;
    assign rom[13'h1a52] = 0;
    assign rom[13'h1a53] = 1;
    assign rom[13'h1a54] = 1;
    assign rom[13'h1a55] = 0;
    assign rom[13'h1a56] = 0;
    assign rom[13'h1a57] = 0;
    assign rom[13'h1a58] = 0;
    assign rom[13'h1a59] = 0;
    assign rom[13'h1a5a] = 0;
    assign rom[13'h1a5b] = 1;
    assign rom[13'h1a5c] = 1;
    assign rom[13'h1a5d] = 0;
    assign rom[13'h1a5e] = 0;
    assign rom[13'h1a5f] = 0;
    assign rom[13'h1a60] = 0;
    assign rom[13'h1a61] = 0;
    assign rom[13'h1a62] = 0;
    assign rom[13'h1a63] = 1;
    assign rom[13'h1a64] = 1;
    assign rom[13'h1a65] = 0;
    assign rom[13'h1a66] = 0;
    assign rom[13'h1a67] = 0;
    assign rom[13'h1a68] = 0;
    assign rom[13'h1a69] = 0;
    assign rom[13'h1a6a] = 0;
    assign rom[13'h1a6b] = 1;
    assign rom[13'h1a6c] = 1;
    assign rom[13'h1a6d] = 0;
    assign rom[13'h1a6e] = 0;
    assign rom[13'h1a6f] = 0;
    assign rom[13'h1a70] = 0;
    assign rom[13'h1a71] = 0;
    assign rom[13'h1a72] = 0;
    assign rom[13'h1a73] = 1;
    assign rom[13'h1a74] = 1;
    assign rom[13'h1a75] = 0;
    assign rom[13'h1a76] = 0;
    assign rom[13'h1a77] = 0;
    assign rom[13'h1a78] = 0;
    assign rom[13'h1a79] = 0;
    assign rom[13'h1a7a] = 0;
    assign rom[13'h1a7b] = 0;
    assign rom[13'h1a7c] = 0;
    assign rom[13'h1a7d] = 0;
    assign rom[13'h1a7e] = 0;
    assign rom[13'h1a7f] = 0;
    assign rom[13'h1a80] = 0;
    assign rom[13'h1a81] = 0;
    assign rom[13'h1a82] = 0;
    assign rom[13'h1a83] = 1;
    assign rom[13'h1a84] = 1;
    assign rom[13'h1a85] = 0;
    assign rom[13'h1a86] = 0;
    assign rom[13'h1a87] = 0;
    assign rom[13'h1a88] = 0;
    assign rom[13'h1a89] = 0;
    assign rom[13'h1a8a] = 0;
    assign rom[13'h1a8b] = 0;
    assign rom[13'h1a8c] = 0;
    assign rom[13'h1a8d] = 0;
    assign rom[13'h1a8e] = 0;
    assign rom[13'h1a8f] = 0;
    assign rom[13'h1a90] = 0;
    assign rom[13'h1a91] = 0;
    assign rom[13'h1a92] = 0;
    assign rom[13'h1a93] = 1;
    assign rom[13'h1a94] = 1;
    assign rom[13'h1a95] = 0;
    assign rom[13'h1a96] = 0;
    assign rom[13'h1a97] = 0;
    assign rom[13'h1a98] = 0;
    assign rom[13'h1a99] = 0;
    assign rom[13'h1a9a] = 0;
    assign rom[13'h1a9b] = 1;
    assign rom[13'h1a9c] = 1;
    assign rom[13'h1a9d] = 0;
    assign rom[13'h1a9e] = 0;
    assign rom[13'h1a9f] = 0;
    assign rom[13'h1aa0] = 0;
    assign rom[13'h1aa1] = 0;
    assign rom[13'h1aa2] = 0;
    assign rom[13'h1aa3] = 1;
    assign rom[13'h1aa4] = 1;
    assign rom[13'h1aa5] = 0;
    assign rom[13'h1aa6] = 0;
    assign rom[13'h1aa7] = 0;
    assign rom[13'h1aa8] = 0;
    assign rom[13'h1aa9] = 0;
    assign rom[13'h1aaa] = 0;
    assign rom[13'h1aab] = 1;
    assign rom[13'h1aac] = 1;
    assign rom[13'h1aad] = 0;
    assign rom[13'h1aae] = 0;
    assign rom[13'h1aaf] = 0;
    assign rom[13'h1ab0] = 0;
    assign rom[13'h1ab1] = 0;
    assign rom[13'h1ab2] = 0;
    assign rom[13'h1ab3] = 1;
    assign rom[13'h1ab4] = 1;
    assign rom[13'h1ab5] = 0;
    assign rom[13'h1ab6] = 0;
    assign rom[13'h1ab7] = 0;
    assign rom[13'h1ab8] = 0;
    assign rom[13'h1ab9] = 1;
    assign rom[13'h1aba] = 1;
    assign rom[13'h1abb] = 1;
    assign rom[13'h1abc] = 0;
    assign rom[13'h1abd] = 0;
    assign rom[13'h1abe] = 0;
    assign rom[13'h1abf] = 0;
    assign rom[13'h1ac0] = 0;
    assign rom[13'h1ac1] = 1;
    assign rom[13'h1ac2] = 1;
    assign rom[13'h1ac3] = 0;
    assign rom[13'h1ac4] = 0;
    assign rom[13'h1ac5] = 0;
    assign rom[13'h1ac6] = 0;
    assign rom[13'h1ac7] = 0;
    assign rom[13'h1ac8] = 0;
    assign rom[13'h1ac9] = 1;
    assign rom[13'h1aca] = 1;
    assign rom[13'h1acb] = 0;
    assign rom[13'h1acc] = 0;
    assign rom[13'h1acd] = 0;
    assign rom[13'h1ace] = 0;
    assign rom[13'h1acf] = 0;
    assign rom[13'h1ad0] = 0;
    assign rom[13'h1ad1] = 1;
    assign rom[13'h1ad2] = 1;
    assign rom[13'h1ad3] = 0;
    assign rom[13'h1ad4] = 0;
    assign rom[13'h1ad5] = 1;
    assign rom[13'h1ad6] = 1;
    assign rom[13'h1ad7] = 0;
    assign rom[13'h1ad8] = 0;
    assign rom[13'h1ad9] = 1;
    assign rom[13'h1ada] = 1;
    assign rom[13'h1adb] = 0;
    assign rom[13'h1adc] = 1;
    assign rom[13'h1add] = 1;
    assign rom[13'h1ade] = 0;
    assign rom[13'h1adf] = 0;
    assign rom[13'h1ae0] = 0;
    assign rom[13'h1ae1] = 1;
    assign rom[13'h1ae2] = 1;
    assign rom[13'h1ae3] = 1;
    assign rom[13'h1ae4] = 1;
    assign rom[13'h1ae5] = 0;
    assign rom[13'h1ae6] = 0;
    assign rom[13'h1ae7] = 0;
    assign rom[13'h1ae8] = 0;
    assign rom[13'h1ae9] = 1;
    assign rom[13'h1aea] = 1;
    assign rom[13'h1aeb] = 0;
    assign rom[13'h1aec] = 1;
    assign rom[13'h1aed] = 1;
    assign rom[13'h1aee] = 0;
    assign rom[13'h1aef] = 0;
    assign rom[13'h1af0] = 0;
    assign rom[13'h1af1] = 1;
    assign rom[13'h1af2] = 1;
    assign rom[13'h1af3] = 0;
    assign rom[13'h1af4] = 0;
    assign rom[13'h1af5] = 1;
    assign rom[13'h1af6] = 1;
    assign rom[13'h1af7] = 0;
    assign rom[13'h1af8] = 0;
    assign rom[13'h1af9] = 0;
    assign rom[13'h1afa] = 0;
    assign rom[13'h1afb] = 0;
    assign rom[13'h1afc] = 0;
    assign rom[13'h1afd] = 0;
    assign rom[13'h1afe] = 0;
    assign rom[13'h1aff] = 0;
    assign rom[13'h1b00] = 0;
    assign rom[13'h1b01] = 0;
    assign rom[13'h1b02] = 1;
    assign rom[13'h1b03] = 1;
    assign rom[13'h1b04] = 0;
    assign rom[13'h1b05] = 0;
    assign rom[13'h1b06] = 0;
    assign rom[13'h1b07] = 0;
    assign rom[13'h1b08] = 0;
    assign rom[13'h1b09] = 0;
    assign rom[13'h1b0a] = 1;
    assign rom[13'h1b0b] = 1;
    assign rom[13'h1b0c] = 0;
    assign rom[13'h1b0d] = 0;
    assign rom[13'h1b0e] = 0;
    assign rom[13'h1b0f] = 0;
    assign rom[13'h1b10] = 0;
    assign rom[13'h1b11] = 0;
    assign rom[13'h1b12] = 1;
    assign rom[13'h1b13] = 1;
    assign rom[13'h1b14] = 0;
    assign rom[13'h1b15] = 0;
    assign rom[13'h1b16] = 0;
    assign rom[13'h1b17] = 0;
    assign rom[13'h1b18] = 0;
    assign rom[13'h1b19] = 0;
    assign rom[13'h1b1a] = 1;
    assign rom[13'h1b1b] = 1;
    assign rom[13'h1b1c] = 0;
    assign rom[13'h1b1d] = 0;
    assign rom[13'h1b1e] = 0;
    assign rom[13'h1b1f] = 0;
    assign rom[13'h1b20] = 0;
    assign rom[13'h1b21] = 0;
    assign rom[13'h1b22] = 1;
    assign rom[13'h1b23] = 1;
    assign rom[13'h1b24] = 0;
    assign rom[13'h1b25] = 0;
    assign rom[13'h1b26] = 0;
    assign rom[13'h1b27] = 0;
    assign rom[13'h1b28] = 0;
    assign rom[13'h1b29] = 0;
    assign rom[13'h1b2a] = 1;
    assign rom[13'h1b2b] = 1;
    assign rom[13'h1b2c] = 0;
    assign rom[13'h1b2d] = 0;
    assign rom[13'h1b2e] = 0;
    assign rom[13'h1b2f] = 0;
    assign rom[13'h1b30] = 0;
    assign rom[13'h1b31] = 0;
    assign rom[13'h1b32] = 0;
    assign rom[13'h1b33] = 1;
    assign rom[13'h1b34] = 1;
    assign rom[13'h1b35] = 1;
    assign rom[13'h1b36] = 0;
    assign rom[13'h1b37] = 0;
    assign rom[13'h1b38] = 0;
    assign rom[13'h1b39] = 0;
    assign rom[13'h1b3a] = 0;
    assign rom[13'h1b3b] = 0;
    assign rom[13'h1b3c] = 0;
    assign rom[13'h1b3d] = 0;
    assign rom[13'h1b3e] = 0;
    assign rom[13'h1b3f] = 0;
    assign rom[13'h1b40] = 0;
    assign rom[13'h1b41] = 0;
    assign rom[13'h1b42] = 0;
    assign rom[13'h1b43] = 0;
    assign rom[13'h1b44] = 0;
    assign rom[13'h1b45] = 0;
    assign rom[13'h1b46] = 0;
    assign rom[13'h1b47] = 0;
    assign rom[13'h1b48] = 0;
    assign rom[13'h1b49] = 0;
    assign rom[13'h1b4a] = 0;
    assign rom[13'h1b4b] = 0;
    assign rom[13'h1b4c] = 0;
    assign rom[13'h1b4d] = 0;
    assign rom[13'h1b4e] = 0;
    assign rom[13'h1b4f] = 0;
    assign rom[13'h1b50] = 1;
    assign rom[13'h1b51] = 1;
    assign rom[13'h1b52] = 0;
    assign rom[13'h1b53] = 0;
    assign rom[13'h1b54] = 1;
    assign rom[13'h1b55] = 1;
    assign rom[13'h1b56] = 0;
    assign rom[13'h1b57] = 0;
    assign rom[13'h1b58] = 1;
    assign rom[13'h1b59] = 1;
    assign rom[13'h1b5a] = 1;
    assign rom[13'h1b5b] = 1;
    assign rom[13'h1b5c] = 1;
    assign rom[13'h1b5d] = 1;
    assign rom[13'h1b5e] = 1;
    assign rom[13'h1b5f] = 0;
    assign rom[13'h1b60] = 1;
    assign rom[13'h1b61] = 1;
    assign rom[13'h1b62] = 0;
    assign rom[13'h1b63] = 1;
    assign rom[13'h1b64] = 0;
    assign rom[13'h1b65] = 1;
    assign rom[13'h1b66] = 1;
    assign rom[13'h1b67] = 0;
    assign rom[13'h1b68] = 1;
    assign rom[13'h1b69] = 1;
    assign rom[13'h1b6a] = 0;
    assign rom[13'h1b6b] = 0;
    assign rom[13'h1b6c] = 0;
    assign rom[13'h1b6d] = 1;
    assign rom[13'h1b6e] = 1;
    assign rom[13'h1b6f] = 0;
    assign rom[13'h1b70] = 1;
    assign rom[13'h1b71] = 1;
    assign rom[13'h1b72] = 0;
    assign rom[13'h1b73] = 0;
    assign rom[13'h1b74] = 0;
    assign rom[13'h1b75] = 1;
    assign rom[13'h1b76] = 1;
    assign rom[13'h1b77] = 0;
    assign rom[13'h1b78] = 0;
    assign rom[13'h1b79] = 0;
    assign rom[13'h1b7a] = 0;
    assign rom[13'h1b7b] = 0;
    assign rom[13'h1b7c] = 0;
    assign rom[13'h1b7d] = 0;
    assign rom[13'h1b7e] = 0;
    assign rom[13'h1b7f] = 0;
    assign rom[13'h1b80] = 0;
    assign rom[13'h1b81] = 0;
    assign rom[13'h1b82] = 0;
    assign rom[13'h1b83] = 0;
    assign rom[13'h1b84] = 0;
    assign rom[13'h1b85] = 0;
    assign rom[13'h1b86] = 0;
    assign rom[13'h1b87] = 0;
    assign rom[13'h1b88] = 0;
    assign rom[13'h1b89] = 0;
    assign rom[13'h1b8a] = 0;
    assign rom[13'h1b8b] = 0;
    assign rom[13'h1b8c] = 0;
    assign rom[13'h1b8d] = 0;
    assign rom[13'h1b8e] = 0;
    assign rom[13'h1b8f] = 0;
    assign rom[13'h1b90] = 0;
    assign rom[13'h1b91] = 1;
    assign rom[13'h1b92] = 1;
    assign rom[13'h1b93] = 1;
    assign rom[13'h1b94] = 1;
    assign rom[13'h1b95] = 1;
    assign rom[13'h1b96] = 0;
    assign rom[13'h1b97] = 0;
    assign rom[13'h1b98] = 0;
    assign rom[13'h1b99] = 1;
    assign rom[13'h1b9a] = 1;
    assign rom[13'h1b9b] = 0;
    assign rom[13'h1b9c] = 0;
    assign rom[13'h1b9d] = 1;
    assign rom[13'h1b9e] = 1;
    assign rom[13'h1b9f] = 0;
    assign rom[13'h1ba0] = 0;
    assign rom[13'h1ba1] = 1;
    assign rom[13'h1ba2] = 1;
    assign rom[13'h1ba3] = 0;
    assign rom[13'h1ba4] = 0;
    assign rom[13'h1ba5] = 1;
    assign rom[13'h1ba6] = 1;
    assign rom[13'h1ba7] = 0;
    assign rom[13'h1ba8] = 0;
    assign rom[13'h1ba9] = 1;
    assign rom[13'h1baa] = 1;
    assign rom[13'h1bab] = 0;
    assign rom[13'h1bac] = 0;
    assign rom[13'h1bad] = 1;
    assign rom[13'h1bae] = 1;
    assign rom[13'h1baf] = 0;
    assign rom[13'h1bb0] = 0;
    assign rom[13'h1bb1] = 1;
    assign rom[13'h1bb2] = 1;
    assign rom[13'h1bb3] = 0;
    assign rom[13'h1bb4] = 0;
    assign rom[13'h1bb5] = 1;
    assign rom[13'h1bb6] = 1;
    assign rom[13'h1bb7] = 0;
    assign rom[13'h1bb8] = 0;
    assign rom[13'h1bb9] = 0;
    assign rom[13'h1bba] = 0;
    assign rom[13'h1bbb] = 0;
    assign rom[13'h1bbc] = 0;
    assign rom[13'h1bbd] = 0;
    assign rom[13'h1bbe] = 0;
    assign rom[13'h1bbf] = 0;
    assign rom[13'h1bc0] = 0;
    assign rom[13'h1bc1] = 0;
    assign rom[13'h1bc2] = 0;
    assign rom[13'h1bc3] = 0;
    assign rom[13'h1bc4] = 0;
    assign rom[13'h1bc5] = 0;
    assign rom[13'h1bc6] = 0;
    assign rom[13'h1bc7] = 0;
    assign rom[13'h1bc8] = 0;
    assign rom[13'h1bc9] = 0;
    assign rom[13'h1bca] = 0;
    assign rom[13'h1bcb] = 0;
    assign rom[13'h1bcc] = 0;
    assign rom[13'h1bcd] = 0;
    assign rom[13'h1bce] = 0;
    assign rom[13'h1bcf] = 0;
    assign rom[13'h1bd0] = 0;
    assign rom[13'h1bd1] = 0;
    assign rom[13'h1bd2] = 1;
    assign rom[13'h1bd3] = 1;
    assign rom[13'h1bd4] = 1;
    assign rom[13'h1bd5] = 1;
    assign rom[13'h1bd6] = 0;
    assign rom[13'h1bd7] = 0;
    assign rom[13'h1bd8] = 0;
    assign rom[13'h1bd9] = 1;
    assign rom[13'h1bda] = 1;
    assign rom[13'h1bdb] = 0;
    assign rom[13'h1bdc] = 0;
    assign rom[13'h1bdd] = 1;
    assign rom[13'h1bde] = 1;
    assign rom[13'h1bdf] = 0;
    assign rom[13'h1be0] = 0;
    assign rom[13'h1be1] = 1;
    assign rom[13'h1be2] = 1;
    assign rom[13'h1be3] = 0;
    assign rom[13'h1be4] = 0;
    assign rom[13'h1be5] = 1;
    assign rom[13'h1be6] = 1;
    assign rom[13'h1be7] = 0;
    assign rom[13'h1be8] = 0;
    assign rom[13'h1be9] = 1;
    assign rom[13'h1bea] = 1;
    assign rom[13'h1beb] = 0;
    assign rom[13'h1bec] = 0;
    assign rom[13'h1bed] = 1;
    assign rom[13'h1bee] = 1;
    assign rom[13'h1bef] = 0;
    assign rom[13'h1bf0] = 0;
    assign rom[13'h1bf1] = 0;
    assign rom[13'h1bf2] = 1;
    assign rom[13'h1bf3] = 1;
    assign rom[13'h1bf4] = 1;
    assign rom[13'h1bf5] = 1;
    assign rom[13'h1bf6] = 0;
    assign rom[13'h1bf7] = 0;
    assign rom[13'h1bf8] = 0;
    assign rom[13'h1bf9] = 0;
    assign rom[13'h1bfa] = 0;
    assign rom[13'h1bfb] = 0;
    assign rom[13'h1bfc] = 0;
    assign rom[13'h1bfd] = 0;
    assign rom[13'h1bfe] = 0;
    assign rom[13'h1bff] = 0;
    assign rom[13'h1c00] = 0;
    assign rom[13'h1c01] = 0;
    assign rom[13'h1c02] = 0;
    assign rom[13'h1c03] = 0;
    assign rom[13'h1c04] = 0;
    assign rom[13'h1c05] = 0;
    assign rom[13'h1c06] = 0;
    assign rom[13'h1c07] = 0;
    assign rom[13'h1c08] = 0;
    assign rom[13'h1c09] = 0;
    assign rom[13'h1c0a] = 0;
    assign rom[13'h1c0b] = 0;
    assign rom[13'h1c0c] = 0;
    assign rom[13'h1c0d] = 0;
    assign rom[13'h1c0e] = 0;
    assign rom[13'h1c0f] = 0;
    assign rom[13'h1c10] = 0;
    assign rom[13'h1c11] = 1;
    assign rom[13'h1c12] = 1;
    assign rom[13'h1c13] = 1;
    assign rom[13'h1c14] = 1;
    assign rom[13'h1c15] = 1;
    assign rom[13'h1c16] = 0;
    assign rom[13'h1c17] = 0;
    assign rom[13'h1c18] = 0;
    assign rom[13'h1c19] = 1;
    assign rom[13'h1c1a] = 1;
    assign rom[13'h1c1b] = 0;
    assign rom[13'h1c1c] = 0;
    assign rom[13'h1c1d] = 1;
    assign rom[13'h1c1e] = 1;
    assign rom[13'h1c1f] = 0;
    assign rom[13'h1c20] = 0;
    assign rom[13'h1c21] = 1;
    assign rom[13'h1c22] = 1;
    assign rom[13'h1c23] = 0;
    assign rom[13'h1c24] = 0;
    assign rom[13'h1c25] = 1;
    assign rom[13'h1c26] = 1;
    assign rom[13'h1c27] = 0;
    assign rom[13'h1c28] = 0;
    assign rom[13'h1c29] = 1;
    assign rom[13'h1c2a] = 1;
    assign rom[13'h1c2b] = 1;
    assign rom[13'h1c2c] = 1;
    assign rom[13'h1c2d] = 1;
    assign rom[13'h1c2e] = 0;
    assign rom[13'h1c2f] = 0;
    assign rom[13'h1c30] = 0;
    assign rom[13'h1c31] = 1;
    assign rom[13'h1c32] = 1;
    assign rom[13'h1c33] = 0;
    assign rom[13'h1c34] = 0;
    assign rom[13'h1c35] = 0;
    assign rom[13'h1c36] = 0;
    assign rom[13'h1c37] = 0;
    assign rom[13'h1c38] = 0;
    assign rom[13'h1c39] = 1;
    assign rom[13'h1c3a] = 1;
    assign rom[13'h1c3b] = 0;
    assign rom[13'h1c3c] = 0;
    assign rom[13'h1c3d] = 0;
    assign rom[13'h1c3e] = 0;
    assign rom[13'h1c3f] = 0;
    assign rom[13'h1c40] = 0;
    assign rom[13'h1c41] = 0;
    assign rom[13'h1c42] = 0;
    assign rom[13'h1c43] = 0;
    assign rom[13'h1c44] = 0;
    assign rom[13'h1c45] = 0;
    assign rom[13'h1c46] = 0;
    assign rom[13'h1c47] = 0;
    assign rom[13'h1c48] = 0;
    assign rom[13'h1c49] = 0;
    assign rom[13'h1c4a] = 0;
    assign rom[13'h1c4b] = 0;
    assign rom[13'h1c4c] = 0;
    assign rom[13'h1c4d] = 0;
    assign rom[13'h1c4e] = 0;
    assign rom[13'h1c4f] = 0;
    assign rom[13'h1c50] = 0;
    assign rom[13'h1c51] = 0;
    assign rom[13'h1c52] = 1;
    assign rom[13'h1c53] = 1;
    assign rom[13'h1c54] = 1;
    assign rom[13'h1c55] = 1;
    assign rom[13'h1c56] = 1;
    assign rom[13'h1c57] = 0;
    assign rom[13'h1c58] = 0;
    assign rom[13'h1c59] = 1;
    assign rom[13'h1c5a] = 1;
    assign rom[13'h1c5b] = 0;
    assign rom[13'h1c5c] = 0;
    assign rom[13'h1c5d] = 1;
    assign rom[13'h1c5e] = 1;
    assign rom[13'h1c5f] = 0;
    assign rom[13'h1c60] = 0;
    assign rom[13'h1c61] = 1;
    assign rom[13'h1c62] = 1;
    assign rom[13'h1c63] = 0;
    assign rom[13'h1c64] = 0;
    assign rom[13'h1c65] = 1;
    assign rom[13'h1c66] = 1;
    assign rom[13'h1c67] = 0;
    assign rom[13'h1c68] = 0;
    assign rom[13'h1c69] = 0;
    assign rom[13'h1c6a] = 1;
    assign rom[13'h1c6b] = 1;
    assign rom[13'h1c6c] = 1;
    assign rom[13'h1c6d] = 1;
    assign rom[13'h1c6e] = 1;
    assign rom[13'h1c6f] = 0;
    assign rom[13'h1c70] = 0;
    assign rom[13'h1c71] = 0;
    assign rom[13'h1c72] = 0;
    assign rom[13'h1c73] = 0;
    assign rom[13'h1c74] = 0;
    assign rom[13'h1c75] = 1;
    assign rom[13'h1c76] = 1;
    assign rom[13'h1c77] = 0;
    assign rom[13'h1c78] = 0;
    assign rom[13'h1c79] = 0;
    assign rom[13'h1c7a] = 0;
    assign rom[13'h1c7b] = 0;
    assign rom[13'h1c7c] = 0;
    assign rom[13'h1c7d] = 1;
    assign rom[13'h1c7e] = 1;
    assign rom[13'h1c7f] = 0;
    assign rom[13'h1c80] = 0;
    assign rom[13'h1c81] = 0;
    assign rom[13'h1c82] = 0;
    assign rom[13'h1c83] = 0;
    assign rom[13'h1c84] = 0;
    assign rom[13'h1c85] = 0;
    assign rom[13'h1c86] = 0;
    assign rom[13'h1c87] = 0;
    assign rom[13'h1c88] = 0;
    assign rom[13'h1c89] = 0;
    assign rom[13'h1c8a] = 0;
    assign rom[13'h1c8b] = 0;
    assign rom[13'h1c8c] = 0;
    assign rom[13'h1c8d] = 0;
    assign rom[13'h1c8e] = 0;
    assign rom[13'h1c8f] = 0;
    assign rom[13'h1c90] = 0;
    assign rom[13'h1c91] = 0;
    assign rom[13'h1c92] = 1;
    assign rom[13'h1c93] = 1;
    assign rom[13'h1c94] = 0;
    assign rom[13'h1c95] = 1;
    assign rom[13'h1c96] = 1;
    assign rom[13'h1c97] = 0;
    assign rom[13'h1c98] = 0;
    assign rom[13'h1c99] = 0;
    assign rom[13'h1c9a] = 1;
    assign rom[13'h1c9b] = 1;
    assign rom[13'h1c9c] = 1;
    assign rom[13'h1c9d] = 0;
    assign rom[13'h1c9e] = 0;
    assign rom[13'h1c9f] = 0;
    assign rom[13'h1ca0] = 0;
    assign rom[13'h1ca1] = 0;
    assign rom[13'h1ca2] = 1;
    assign rom[13'h1ca3] = 1;
    assign rom[13'h1ca4] = 0;
    assign rom[13'h1ca5] = 0;
    assign rom[13'h1ca6] = 0;
    assign rom[13'h1ca7] = 0;
    assign rom[13'h1ca8] = 0;
    assign rom[13'h1ca9] = 0;
    assign rom[13'h1caa] = 1;
    assign rom[13'h1cab] = 1;
    assign rom[13'h1cac] = 0;
    assign rom[13'h1cad] = 0;
    assign rom[13'h1cae] = 0;
    assign rom[13'h1caf] = 0;
    assign rom[13'h1cb0] = 0;
    assign rom[13'h1cb1] = 0;
    assign rom[13'h1cb2] = 1;
    assign rom[13'h1cb3] = 1;
    assign rom[13'h1cb4] = 0;
    assign rom[13'h1cb5] = 0;
    assign rom[13'h1cb6] = 0;
    assign rom[13'h1cb7] = 0;
    assign rom[13'h1cb8] = 0;
    assign rom[13'h1cb9] = 0;
    assign rom[13'h1cba] = 0;
    assign rom[13'h1cbb] = 0;
    assign rom[13'h1cbc] = 0;
    assign rom[13'h1cbd] = 0;
    assign rom[13'h1cbe] = 0;
    assign rom[13'h1cbf] = 0;
    assign rom[13'h1cc0] = 0;
    assign rom[13'h1cc1] = 0;
    assign rom[13'h1cc2] = 0;
    assign rom[13'h1cc3] = 0;
    assign rom[13'h1cc4] = 0;
    assign rom[13'h1cc5] = 0;
    assign rom[13'h1cc6] = 0;
    assign rom[13'h1cc7] = 0;
    assign rom[13'h1cc8] = 0;
    assign rom[13'h1cc9] = 0;
    assign rom[13'h1cca] = 0;
    assign rom[13'h1ccb] = 0;
    assign rom[13'h1ccc] = 0;
    assign rom[13'h1ccd] = 0;
    assign rom[13'h1cce] = 0;
    assign rom[13'h1ccf] = 0;
    assign rom[13'h1cd0] = 0;
    assign rom[13'h1cd1] = 0;
    assign rom[13'h1cd2] = 1;
    assign rom[13'h1cd3] = 1;
    assign rom[13'h1cd4] = 1;
    assign rom[13'h1cd5] = 1;
    assign rom[13'h1cd6] = 1;
    assign rom[13'h1cd7] = 0;
    assign rom[13'h1cd8] = 0;
    assign rom[13'h1cd9] = 1;
    assign rom[13'h1cda] = 1;
    assign rom[13'h1cdb] = 0;
    assign rom[13'h1cdc] = 0;
    assign rom[13'h1cdd] = 0;
    assign rom[13'h1cde] = 0;
    assign rom[13'h1cdf] = 0;
    assign rom[13'h1ce0] = 0;
    assign rom[13'h1ce1] = 0;
    assign rom[13'h1ce2] = 1;
    assign rom[13'h1ce3] = 1;
    assign rom[13'h1ce4] = 1;
    assign rom[13'h1ce5] = 1;
    assign rom[13'h1ce6] = 0;
    assign rom[13'h1ce7] = 0;
    assign rom[13'h1ce8] = 0;
    assign rom[13'h1ce9] = 0;
    assign rom[13'h1cea] = 0;
    assign rom[13'h1ceb] = 0;
    assign rom[13'h1cec] = 0;
    assign rom[13'h1ced] = 1;
    assign rom[13'h1cee] = 1;
    assign rom[13'h1cef] = 0;
    assign rom[13'h1cf0] = 0;
    assign rom[13'h1cf1] = 1;
    assign rom[13'h1cf2] = 1;
    assign rom[13'h1cf3] = 1;
    assign rom[13'h1cf4] = 1;
    assign rom[13'h1cf5] = 1;
    assign rom[13'h1cf6] = 0;
    assign rom[13'h1cf7] = 0;
    assign rom[13'h1cf8] = 0;
    assign rom[13'h1cf9] = 0;
    assign rom[13'h1cfa] = 0;
    assign rom[13'h1cfb] = 0;
    assign rom[13'h1cfc] = 0;
    assign rom[13'h1cfd] = 0;
    assign rom[13'h1cfe] = 0;
    assign rom[13'h1cff] = 0;
    assign rom[13'h1d00] = 0;
    assign rom[13'h1d01] = 0;
    assign rom[13'h1d02] = 0;
    assign rom[13'h1d03] = 1;
    assign rom[13'h1d04] = 1;
    assign rom[13'h1d05] = 0;
    assign rom[13'h1d06] = 0;
    assign rom[13'h1d07] = 0;
    assign rom[13'h1d08] = 0;
    assign rom[13'h1d09] = 0;
    assign rom[13'h1d0a] = 0;
    assign rom[13'h1d0b] = 1;
    assign rom[13'h1d0c] = 1;
    assign rom[13'h1d0d] = 0;
    assign rom[13'h1d0e] = 0;
    assign rom[13'h1d0f] = 0;
    assign rom[13'h1d10] = 0;
    assign rom[13'h1d11] = 0;
    assign rom[13'h1d12] = 1;
    assign rom[13'h1d13] = 1;
    assign rom[13'h1d14] = 1;
    assign rom[13'h1d15] = 1;
    assign rom[13'h1d16] = 0;
    assign rom[13'h1d17] = 0;
    assign rom[13'h1d18] = 0;
    assign rom[13'h1d19] = 0;
    assign rom[13'h1d1a] = 0;
    assign rom[13'h1d1b] = 1;
    assign rom[13'h1d1c] = 1;
    assign rom[13'h1d1d] = 0;
    assign rom[13'h1d1e] = 0;
    assign rom[13'h1d1f] = 0;
    assign rom[13'h1d20] = 0;
    assign rom[13'h1d21] = 0;
    assign rom[13'h1d22] = 0;
    assign rom[13'h1d23] = 1;
    assign rom[13'h1d24] = 1;
    assign rom[13'h1d25] = 0;
    assign rom[13'h1d26] = 0;
    assign rom[13'h1d27] = 0;
    assign rom[13'h1d28] = 0;
    assign rom[13'h1d29] = 0;
    assign rom[13'h1d2a] = 0;
    assign rom[13'h1d2b] = 1;
    assign rom[13'h1d2c] = 1;
    assign rom[13'h1d2d] = 0;
    assign rom[13'h1d2e] = 0;
    assign rom[13'h1d2f] = 0;
    assign rom[13'h1d30] = 0;
    assign rom[13'h1d31] = 0;
    assign rom[13'h1d32] = 0;
    assign rom[13'h1d33] = 0;
    assign rom[13'h1d34] = 1;
    assign rom[13'h1d35] = 1;
    assign rom[13'h1d36] = 0;
    assign rom[13'h1d37] = 0;
    assign rom[13'h1d38] = 0;
    assign rom[13'h1d39] = 0;
    assign rom[13'h1d3a] = 0;
    assign rom[13'h1d3b] = 0;
    assign rom[13'h1d3c] = 0;
    assign rom[13'h1d3d] = 0;
    assign rom[13'h1d3e] = 0;
    assign rom[13'h1d3f] = 0;
    assign rom[13'h1d40] = 0;
    assign rom[13'h1d41] = 0;
    assign rom[13'h1d42] = 0;
    assign rom[13'h1d43] = 0;
    assign rom[13'h1d44] = 0;
    assign rom[13'h1d45] = 0;
    assign rom[13'h1d46] = 0;
    assign rom[13'h1d47] = 0;
    assign rom[13'h1d48] = 0;
    assign rom[13'h1d49] = 0;
    assign rom[13'h1d4a] = 0;
    assign rom[13'h1d4b] = 0;
    assign rom[13'h1d4c] = 0;
    assign rom[13'h1d4d] = 0;
    assign rom[13'h1d4e] = 0;
    assign rom[13'h1d4f] = 0;
    assign rom[13'h1d50] = 0;
    assign rom[13'h1d51] = 1;
    assign rom[13'h1d52] = 1;
    assign rom[13'h1d53] = 0;
    assign rom[13'h1d54] = 0;
    assign rom[13'h1d55] = 1;
    assign rom[13'h1d56] = 1;
    assign rom[13'h1d57] = 0;
    assign rom[13'h1d58] = 0;
    assign rom[13'h1d59] = 1;
    assign rom[13'h1d5a] = 1;
    assign rom[13'h1d5b] = 0;
    assign rom[13'h1d5c] = 0;
    assign rom[13'h1d5d] = 1;
    assign rom[13'h1d5e] = 1;
    assign rom[13'h1d5f] = 0;
    assign rom[13'h1d60] = 0;
    assign rom[13'h1d61] = 1;
    assign rom[13'h1d62] = 1;
    assign rom[13'h1d63] = 0;
    assign rom[13'h1d64] = 0;
    assign rom[13'h1d65] = 1;
    assign rom[13'h1d66] = 1;
    assign rom[13'h1d67] = 0;
    assign rom[13'h1d68] = 0;
    assign rom[13'h1d69] = 1;
    assign rom[13'h1d6a] = 1;
    assign rom[13'h1d6b] = 0;
    assign rom[13'h1d6c] = 0;
    assign rom[13'h1d6d] = 1;
    assign rom[13'h1d6e] = 1;
    assign rom[13'h1d6f] = 0;
    assign rom[13'h1d70] = 0;
    assign rom[13'h1d71] = 0;
    assign rom[13'h1d72] = 1;
    assign rom[13'h1d73] = 1;
    assign rom[13'h1d74] = 1;
    assign rom[13'h1d75] = 1;
    assign rom[13'h1d76] = 0;
    assign rom[13'h1d77] = 0;
    assign rom[13'h1d78] = 0;
    assign rom[13'h1d79] = 0;
    assign rom[13'h1d7a] = 0;
    assign rom[13'h1d7b] = 0;
    assign rom[13'h1d7c] = 0;
    assign rom[13'h1d7d] = 0;
    assign rom[13'h1d7e] = 0;
    assign rom[13'h1d7f] = 0;
    assign rom[13'h1d80] = 0;
    assign rom[13'h1d81] = 0;
    assign rom[13'h1d82] = 0;
    assign rom[13'h1d83] = 0;
    assign rom[13'h1d84] = 0;
    assign rom[13'h1d85] = 0;
    assign rom[13'h1d86] = 0;
    assign rom[13'h1d87] = 0;
    assign rom[13'h1d88] = 0;
    assign rom[13'h1d89] = 0;
    assign rom[13'h1d8a] = 0;
    assign rom[13'h1d8b] = 0;
    assign rom[13'h1d8c] = 0;
    assign rom[13'h1d8d] = 0;
    assign rom[13'h1d8e] = 0;
    assign rom[13'h1d8f] = 0;
    assign rom[13'h1d90] = 0;
    assign rom[13'h1d91] = 1;
    assign rom[13'h1d92] = 1;
    assign rom[13'h1d93] = 0;
    assign rom[13'h1d94] = 0;
    assign rom[13'h1d95] = 1;
    assign rom[13'h1d96] = 1;
    assign rom[13'h1d97] = 0;
    assign rom[13'h1d98] = 0;
    assign rom[13'h1d99] = 1;
    assign rom[13'h1d9a] = 1;
    assign rom[13'h1d9b] = 0;
    assign rom[13'h1d9c] = 0;
    assign rom[13'h1d9d] = 1;
    assign rom[13'h1d9e] = 1;
    assign rom[13'h1d9f] = 0;
    assign rom[13'h1da0] = 0;
    assign rom[13'h1da1] = 1;
    assign rom[13'h1da2] = 1;
    assign rom[13'h1da3] = 0;
    assign rom[13'h1da4] = 0;
    assign rom[13'h1da5] = 1;
    assign rom[13'h1da6] = 1;
    assign rom[13'h1da7] = 0;
    assign rom[13'h1da8] = 0;
    assign rom[13'h1da9] = 0;
    assign rom[13'h1daa] = 1;
    assign rom[13'h1dab] = 1;
    assign rom[13'h1dac] = 1;
    assign rom[13'h1dad] = 1;
    assign rom[13'h1dae] = 0;
    assign rom[13'h1daf] = 0;
    assign rom[13'h1db0] = 0;
    assign rom[13'h1db1] = 0;
    assign rom[13'h1db2] = 0;
    assign rom[13'h1db3] = 1;
    assign rom[13'h1db4] = 1;
    assign rom[13'h1db5] = 0;
    assign rom[13'h1db6] = 0;
    assign rom[13'h1db7] = 0;
    assign rom[13'h1db8] = 0;
    assign rom[13'h1db9] = 0;
    assign rom[13'h1dba] = 0;
    assign rom[13'h1dbb] = 0;
    assign rom[13'h1dbc] = 0;
    assign rom[13'h1dbd] = 0;
    assign rom[13'h1dbe] = 0;
    assign rom[13'h1dbf] = 0;
    assign rom[13'h1dc0] = 0;
    assign rom[13'h1dc1] = 0;
    assign rom[13'h1dc2] = 0;
    assign rom[13'h1dc3] = 0;
    assign rom[13'h1dc4] = 0;
    assign rom[13'h1dc5] = 0;
    assign rom[13'h1dc6] = 0;
    assign rom[13'h1dc7] = 0;
    assign rom[13'h1dc8] = 0;
    assign rom[13'h1dc9] = 0;
    assign rom[13'h1dca] = 0;
    assign rom[13'h1dcb] = 0;
    assign rom[13'h1dcc] = 0;
    assign rom[13'h1dcd] = 0;
    assign rom[13'h1dce] = 0;
    assign rom[13'h1dcf] = 0;
    assign rom[13'h1dd0] = 1;
    assign rom[13'h1dd1] = 1;
    assign rom[13'h1dd2] = 0;
    assign rom[13'h1dd3] = 0;
    assign rom[13'h1dd4] = 0;
    assign rom[13'h1dd5] = 1;
    assign rom[13'h1dd6] = 1;
    assign rom[13'h1dd7] = 0;
    assign rom[13'h1dd8] = 1;
    assign rom[13'h1dd9] = 1;
    assign rom[13'h1dda] = 0;
    assign rom[13'h1ddb] = 1;
    assign rom[13'h1ddc] = 0;
    assign rom[13'h1ddd] = 1;
    assign rom[13'h1dde] = 1;
    assign rom[13'h1ddf] = 0;
    assign rom[13'h1de0] = 1;
    assign rom[13'h1de1] = 1;
    assign rom[13'h1de2] = 0;
    assign rom[13'h1de3] = 1;
    assign rom[13'h1de4] = 0;
    assign rom[13'h1de5] = 1;
    assign rom[13'h1de6] = 1;
    assign rom[13'h1de7] = 0;
    assign rom[13'h1de8] = 0;
    assign rom[13'h1de9] = 1;
    assign rom[13'h1dea] = 1;
    assign rom[13'h1deb] = 1;
    assign rom[13'h1dec] = 1;
    assign rom[13'h1ded] = 1;
    assign rom[13'h1dee] = 0;
    assign rom[13'h1def] = 0;
    assign rom[13'h1df0] = 0;
    assign rom[13'h1df1] = 0;
    assign rom[13'h1df2] = 1;
    assign rom[13'h1df3] = 0;
    assign rom[13'h1df4] = 1;
    assign rom[13'h1df5] = 0;
    assign rom[13'h1df6] = 0;
    assign rom[13'h1df7] = 0;
    assign rom[13'h1df8] = 0;
    assign rom[13'h1df9] = 0;
    assign rom[13'h1dfa] = 0;
    assign rom[13'h1dfb] = 0;
    assign rom[13'h1dfc] = 0;
    assign rom[13'h1dfd] = 0;
    assign rom[13'h1dfe] = 0;
    assign rom[13'h1dff] = 0;
    assign rom[13'h1e00] = 0;
    assign rom[13'h1e01] = 0;
    assign rom[13'h1e02] = 0;
    assign rom[13'h1e03] = 0;
    assign rom[13'h1e04] = 0;
    assign rom[13'h1e05] = 0;
    assign rom[13'h1e06] = 0;
    assign rom[13'h1e07] = 0;
    assign rom[13'h1e08] = 0;
    assign rom[13'h1e09] = 0;
    assign rom[13'h1e0a] = 0;
    assign rom[13'h1e0b] = 0;
    assign rom[13'h1e0c] = 0;
    assign rom[13'h1e0d] = 0;
    assign rom[13'h1e0e] = 0;
    assign rom[13'h1e0f] = 0;
    assign rom[13'h1e10] = 0;
    assign rom[13'h1e11] = 1;
    assign rom[13'h1e12] = 1;
    assign rom[13'h1e13] = 0;
    assign rom[13'h1e14] = 0;
    assign rom[13'h1e15] = 1;
    assign rom[13'h1e16] = 1;
    assign rom[13'h1e17] = 0;
    assign rom[13'h1e18] = 0;
    assign rom[13'h1e19] = 0;
    assign rom[13'h1e1a] = 1;
    assign rom[13'h1e1b] = 1;
    assign rom[13'h1e1c] = 1;
    assign rom[13'h1e1d] = 1;
    assign rom[13'h1e1e] = 0;
    assign rom[13'h1e1f] = 0;
    assign rom[13'h1e20] = 0;
    assign rom[13'h1e21] = 0;
    assign rom[13'h1e22] = 0;
    assign rom[13'h1e23] = 1;
    assign rom[13'h1e24] = 1;
    assign rom[13'h1e25] = 0;
    assign rom[13'h1e26] = 0;
    assign rom[13'h1e27] = 0;
    assign rom[13'h1e28] = 0;
    assign rom[13'h1e29] = 0;
    assign rom[13'h1e2a] = 1;
    assign rom[13'h1e2b] = 1;
    assign rom[13'h1e2c] = 1;
    assign rom[13'h1e2d] = 1;
    assign rom[13'h1e2e] = 0;
    assign rom[13'h1e2f] = 0;
    assign rom[13'h1e30] = 0;
    assign rom[13'h1e31] = 1;
    assign rom[13'h1e32] = 1;
    assign rom[13'h1e33] = 0;
    assign rom[13'h1e34] = 0;
    assign rom[13'h1e35] = 1;
    assign rom[13'h1e36] = 1;
    assign rom[13'h1e37] = 0;
    assign rom[13'h1e38] = 0;
    assign rom[13'h1e39] = 0;
    assign rom[13'h1e3a] = 0;
    assign rom[13'h1e3b] = 0;
    assign rom[13'h1e3c] = 0;
    assign rom[13'h1e3d] = 0;
    assign rom[13'h1e3e] = 0;
    assign rom[13'h1e3f] = 0;
    assign rom[13'h1e40] = 0;
    assign rom[13'h1e41] = 0;
    assign rom[13'h1e42] = 0;
    assign rom[13'h1e43] = 0;
    assign rom[13'h1e44] = 0;
    assign rom[13'h1e45] = 0;
    assign rom[13'h1e46] = 0;
    assign rom[13'h1e47] = 0;
    assign rom[13'h1e48] = 0;
    assign rom[13'h1e49] = 0;
    assign rom[13'h1e4a] = 0;
    assign rom[13'h1e4b] = 0;
    assign rom[13'h1e4c] = 0;
    assign rom[13'h1e4d] = 0;
    assign rom[13'h1e4e] = 0;
    assign rom[13'h1e4f] = 0;
    assign rom[13'h1e50] = 0;
    assign rom[13'h1e51] = 1;
    assign rom[13'h1e52] = 1;
    assign rom[13'h1e53] = 0;
    assign rom[13'h1e54] = 0;
    assign rom[13'h1e55] = 1;
    assign rom[13'h1e56] = 1;
    assign rom[13'h1e57] = 0;
    assign rom[13'h1e58] = 0;
    assign rom[13'h1e59] = 1;
    assign rom[13'h1e5a] = 1;
    assign rom[13'h1e5b] = 0;
    assign rom[13'h1e5c] = 0;
    assign rom[13'h1e5d] = 1;
    assign rom[13'h1e5e] = 1;
    assign rom[13'h1e5f] = 0;
    assign rom[13'h1e60] = 0;
    assign rom[13'h1e61] = 1;
    assign rom[13'h1e62] = 1;
    assign rom[13'h1e63] = 0;
    assign rom[13'h1e64] = 0;
    assign rom[13'h1e65] = 1;
    assign rom[13'h1e66] = 1;
    assign rom[13'h1e67] = 0;
    assign rom[13'h1e68] = 0;
    assign rom[13'h1e69] = 0;
    assign rom[13'h1e6a] = 1;
    assign rom[13'h1e6b] = 1;
    assign rom[13'h1e6c] = 1;
    assign rom[13'h1e6d] = 1;
    assign rom[13'h1e6e] = 1;
    assign rom[13'h1e6f] = 0;
    assign rom[13'h1e70] = 0;
    assign rom[13'h1e71] = 0;
    assign rom[13'h1e72] = 0;
    assign rom[13'h1e73] = 0;
    assign rom[13'h1e74] = 0;
    assign rom[13'h1e75] = 1;
    assign rom[13'h1e76] = 1;
    assign rom[13'h1e77] = 0;
    assign rom[13'h1e78] = 0;
    assign rom[13'h1e79] = 1;
    assign rom[13'h1e7a] = 1;
    assign rom[13'h1e7b] = 1;
    assign rom[13'h1e7c] = 1;
    assign rom[13'h1e7d] = 1;
    assign rom[13'h1e7e] = 0;
    assign rom[13'h1e7f] = 0;
    assign rom[13'h1e80] = 0;
    assign rom[13'h1e81] = 0;
    assign rom[13'h1e82] = 0;
    assign rom[13'h1e83] = 0;
    assign rom[13'h1e84] = 0;
    assign rom[13'h1e85] = 0;
    assign rom[13'h1e86] = 0;
    assign rom[13'h1e87] = 0;
    assign rom[13'h1e88] = 0;
    assign rom[13'h1e89] = 0;
    assign rom[13'h1e8a] = 0;
    assign rom[13'h1e8b] = 0;
    assign rom[13'h1e8c] = 0;
    assign rom[13'h1e8d] = 0;
    assign rom[13'h1e8e] = 0;
    assign rom[13'h1e8f] = 0;
    assign rom[13'h1e90] = 0;
    assign rom[13'h1e91] = 1;
    assign rom[13'h1e92] = 1;
    assign rom[13'h1e93] = 1;
    assign rom[13'h1e94] = 1;
    assign rom[13'h1e95] = 1;
    assign rom[13'h1e96] = 1;
    assign rom[13'h1e97] = 0;
    assign rom[13'h1e98] = 0;
    assign rom[13'h1e99] = 0;
    assign rom[13'h1e9a] = 0;
    assign rom[13'h1e9b] = 0;
    assign rom[13'h1e9c] = 1;
    assign rom[13'h1e9d] = 1;
    assign rom[13'h1e9e] = 0;
    assign rom[13'h1e9f] = 0;
    assign rom[13'h1ea0] = 0;
    assign rom[13'h1ea1] = 0;
    assign rom[13'h1ea2] = 0;
    assign rom[13'h1ea3] = 1;
    assign rom[13'h1ea4] = 1;
    assign rom[13'h1ea5] = 0;
    assign rom[13'h1ea6] = 0;
    assign rom[13'h1ea7] = 0;
    assign rom[13'h1ea8] = 0;
    assign rom[13'h1ea9] = 0;
    assign rom[13'h1eaa] = 1;
    assign rom[13'h1eab] = 1;
    assign rom[13'h1eac] = 0;
    assign rom[13'h1ead] = 0;
    assign rom[13'h1eae] = 0;
    assign rom[13'h1eaf] = 0;
    assign rom[13'h1eb0] = 0;
    assign rom[13'h1eb1] = 1;
    assign rom[13'h1eb2] = 1;
    assign rom[13'h1eb3] = 1;
    assign rom[13'h1eb4] = 1;
    assign rom[13'h1eb5] = 1;
    assign rom[13'h1eb6] = 1;
    assign rom[13'h1eb7] = 0;
    assign rom[13'h1eb8] = 0;
    assign rom[13'h1eb9] = 0;
    assign rom[13'h1eba] = 0;
    assign rom[13'h1ebb] = 0;
    assign rom[13'h1ebc] = 0;
    assign rom[13'h1ebd] = 0;
    assign rom[13'h1ebe] = 0;
    assign rom[13'h1ebf] = 0;
    assign rom[13'h1ec0] = 0;
    assign rom[13'h1ec1] = 0;
    assign rom[13'h1ec2] = 0;
    assign rom[13'h1ec3] = 1;
    assign rom[13'h1ec4] = 1;
    assign rom[13'h1ec5] = 1;
    assign rom[13'h1ec6] = 0;
    assign rom[13'h1ec7] = 0;
    assign rom[13'h1ec8] = 0;
    assign rom[13'h1ec9] = 0;
    assign rom[13'h1eca] = 1;
    assign rom[13'h1ecb] = 1;
    assign rom[13'h1ecc] = 0;
    assign rom[13'h1ecd] = 0;
    assign rom[13'h1ece] = 0;
    assign rom[13'h1ecf] = 0;
    assign rom[13'h1ed0] = 0;
    assign rom[13'h1ed1] = 0;
    assign rom[13'h1ed2] = 1;
    assign rom[13'h1ed3] = 1;
    assign rom[13'h1ed4] = 0;
    assign rom[13'h1ed5] = 0;
    assign rom[13'h1ed6] = 0;
    assign rom[13'h1ed7] = 0;
    assign rom[13'h1ed8] = 0;
    assign rom[13'h1ed9] = 1;
    assign rom[13'h1eda] = 1;
    assign rom[13'h1edb] = 0;
    assign rom[13'h1edc] = 0;
    assign rom[13'h1edd] = 0;
    assign rom[13'h1ede] = 0;
    assign rom[13'h1edf] = 0;
    assign rom[13'h1ee0] = 0;
    assign rom[13'h1ee1] = 0;
    assign rom[13'h1ee2] = 1;
    assign rom[13'h1ee3] = 1;
    assign rom[13'h1ee4] = 0;
    assign rom[13'h1ee5] = 0;
    assign rom[13'h1ee6] = 0;
    assign rom[13'h1ee7] = 0;
    assign rom[13'h1ee8] = 0;
    assign rom[13'h1ee9] = 0;
    assign rom[13'h1eea] = 1;
    assign rom[13'h1eeb] = 1;
    assign rom[13'h1eec] = 0;
    assign rom[13'h1eed] = 0;
    assign rom[13'h1eee] = 0;
    assign rom[13'h1eef] = 0;
    assign rom[13'h1ef0] = 0;
    assign rom[13'h1ef1] = 0;
    assign rom[13'h1ef2] = 0;
    assign rom[13'h1ef3] = 1;
    assign rom[13'h1ef4] = 1;
    assign rom[13'h1ef5] = 1;
    assign rom[13'h1ef6] = 0;
    assign rom[13'h1ef7] = 0;
    assign rom[13'h1ef8] = 0;
    assign rom[13'h1ef9] = 0;
    assign rom[13'h1efa] = 0;
    assign rom[13'h1efb] = 0;
    assign rom[13'h1efc] = 0;
    assign rom[13'h1efd] = 0;
    assign rom[13'h1efe] = 0;
    assign rom[13'h1eff] = 0;
    assign rom[13'h1f00] = 0;
    assign rom[13'h1f01] = 0;
    assign rom[13'h1f02] = 0;
    assign rom[13'h1f03] = 1;
    assign rom[13'h1f04] = 1;
    assign rom[13'h1f05] = 0;
    assign rom[13'h1f06] = 0;
    assign rom[13'h1f07] = 0;
    assign rom[13'h1f08] = 0;
    assign rom[13'h1f09] = 0;
    assign rom[13'h1f0a] = 0;
    assign rom[13'h1f0b] = 1;
    assign rom[13'h1f0c] = 1;
    assign rom[13'h1f0d] = 0;
    assign rom[13'h1f0e] = 0;
    assign rom[13'h1f0f] = 0;
    assign rom[13'h1f10] = 0;
    assign rom[13'h1f11] = 0;
    assign rom[13'h1f12] = 0;
    assign rom[13'h1f13] = 1;
    assign rom[13'h1f14] = 1;
    assign rom[13'h1f15] = 0;
    assign rom[13'h1f16] = 0;
    assign rom[13'h1f17] = 0;
    assign rom[13'h1f18] = 0;
    assign rom[13'h1f19] = 0;
    assign rom[13'h1f1a] = 0;
    assign rom[13'h1f1b] = 1;
    assign rom[13'h1f1c] = 1;
    assign rom[13'h1f1d] = 0;
    assign rom[13'h1f1e] = 0;
    assign rom[13'h1f1f] = 0;
    assign rom[13'h1f20] = 0;
    assign rom[13'h1f21] = 0;
    assign rom[13'h1f22] = 0;
    assign rom[13'h1f23] = 1;
    assign rom[13'h1f24] = 1;
    assign rom[13'h1f25] = 0;
    assign rom[13'h1f26] = 0;
    assign rom[13'h1f27] = 0;
    assign rom[13'h1f28] = 0;
    assign rom[13'h1f29] = 0;
    assign rom[13'h1f2a] = 0;
    assign rom[13'h1f2b] = 1;
    assign rom[13'h1f2c] = 1;
    assign rom[13'h1f2d] = 0;
    assign rom[13'h1f2e] = 0;
    assign rom[13'h1f2f] = 0;
    assign rom[13'h1f30] = 0;
    assign rom[13'h1f31] = 0;
    assign rom[13'h1f32] = 0;
    assign rom[13'h1f33] = 1;
    assign rom[13'h1f34] = 1;
    assign rom[13'h1f35] = 0;
    assign rom[13'h1f36] = 0;
    assign rom[13'h1f37] = 0;
    assign rom[13'h1f38] = 0;
    assign rom[13'h1f39] = 0;
    assign rom[13'h1f3a] = 0;
    assign rom[13'h1f3b] = 0;
    assign rom[13'h1f3c] = 0;
    assign rom[13'h1f3d] = 0;
    assign rom[13'h1f3e] = 0;
    assign rom[13'h1f3f] = 0;
    assign rom[13'h1f40] = 0;
    assign rom[13'h1f41] = 0;
    assign rom[13'h1f42] = 1;
    assign rom[13'h1f43] = 1;
    assign rom[13'h1f44] = 1;
    assign rom[13'h1f45] = 0;
    assign rom[13'h1f46] = 0;
    assign rom[13'h1f47] = 0;
    assign rom[13'h1f48] = 0;
    assign rom[13'h1f49] = 0;
    assign rom[13'h1f4a] = 0;
    assign rom[13'h1f4b] = 0;
    assign rom[13'h1f4c] = 1;
    assign rom[13'h1f4d] = 1;
    assign rom[13'h1f4e] = 0;
    assign rom[13'h1f4f] = 0;
    assign rom[13'h1f50] = 0;
    assign rom[13'h1f51] = 0;
    assign rom[13'h1f52] = 0;
    assign rom[13'h1f53] = 0;
    assign rom[13'h1f54] = 1;
    assign rom[13'h1f55] = 1;
    assign rom[13'h1f56] = 0;
    assign rom[13'h1f57] = 0;
    assign rom[13'h1f58] = 0;
    assign rom[13'h1f59] = 0;
    assign rom[13'h1f5a] = 0;
    assign rom[13'h1f5b] = 0;
    assign rom[13'h1f5c] = 0;
    assign rom[13'h1f5d] = 1;
    assign rom[13'h1f5e] = 1;
    assign rom[13'h1f5f] = 0;
    assign rom[13'h1f60] = 0;
    assign rom[13'h1f61] = 0;
    assign rom[13'h1f62] = 0;
    assign rom[13'h1f63] = 0;
    assign rom[13'h1f64] = 1;
    assign rom[13'h1f65] = 1;
    assign rom[13'h1f66] = 0;
    assign rom[13'h1f67] = 0;
    assign rom[13'h1f68] = 0;
    assign rom[13'h1f69] = 0;
    assign rom[13'h1f6a] = 0;
    assign rom[13'h1f6b] = 0;
    assign rom[13'h1f6c] = 1;
    assign rom[13'h1f6d] = 1;
    assign rom[13'h1f6e] = 0;
    assign rom[13'h1f6f] = 0;
    assign rom[13'h1f70] = 0;
    assign rom[13'h1f71] = 0;
    assign rom[13'h1f72] = 1;
    assign rom[13'h1f73] = 1;
    assign rom[13'h1f74] = 1;
    assign rom[13'h1f75] = 0;
    assign rom[13'h1f76] = 0;
    assign rom[13'h1f77] = 0;
    assign rom[13'h1f78] = 0;
    assign rom[13'h1f79] = 0;
    assign rom[13'h1f7a] = 0;
    assign rom[13'h1f7b] = 0;
    assign rom[13'h1f7c] = 0;
    assign rom[13'h1f7d] = 0;
    assign rom[13'h1f7e] = 0;
    assign rom[13'h1f7f] = 0;
    assign rom[13'h1f80] = 0;
    assign rom[13'h1f81] = 0;
    assign rom[13'h1f82] = 0;
    assign rom[13'h1f83] = 0;
    assign rom[13'h1f84] = 0;
    assign rom[13'h1f85] = 0;
    assign rom[13'h1f86] = 0;
    assign rom[13'h1f87] = 0;
    assign rom[13'h1f88] = 0;
    assign rom[13'h1f89] = 0;
    assign rom[13'h1f8a] = 1;
    assign rom[13'h1f8b] = 1;
    assign rom[13'h1f8c] = 0;
    assign rom[13'h1f8d] = 0;
    assign rom[13'h1f8e] = 1;
    assign rom[13'h1f8f] = 0;
    assign rom[13'h1f90] = 0;
    assign rom[13'h1f91] = 1;
    assign rom[13'h1f92] = 0;
    assign rom[13'h1f93] = 0;
    assign rom[13'h1f94] = 1;
    assign rom[13'h1f95] = 1;
    assign rom[13'h1f96] = 0;
    assign rom[13'h1f97] = 0;
    assign rom[13'h1f98] = 0;
    assign rom[13'h1f99] = 0;
    assign rom[13'h1f9a] = 0;
    assign rom[13'h1f9b] = 0;
    assign rom[13'h1f9c] = 0;
    assign rom[13'h1f9d] = 0;
    assign rom[13'h1f9e] = 0;
    assign rom[13'h1f9f] = 0;
    assign rom[13'h1fa0] = 0;
    assign rom[13'h1fa1] = 0;
    assign rom[13'h1fa2] = 0;
    assign rom[13'h1fa3] = 0;
    assign rom[13'h1fa4] = 0;
    assign rom[13'h1fa5] = 0;
    assign rom[13'h1fa6] = 0;
    assign rom[13'h1fa7] = 0;
    assign rom[13'h1fa8] = 0;
    assign rom[13'h1fa9] = 0;
    assign rom[13'h1faa] = 0;
    assign rom[13'h1fab] = 0;
    assign rom[13'h1fac] = 0;
    assign rom[13'h1fad] = 0;
    assign rom[13'h1fae] = 0;
    assign rom[13'h1faf] = 0;
    assign rom[13'h1fb0] = 0;
    assign rom[13'h1fb1] = 0;
    assign rom[13'h1fb2] = 0;
    assign rom[13'h1fb3] = 0;
    assign rom[13'h1fb4] = 0;
    assign rom[13'h1fb5] = 0;
    assign rom[13'h1fb6] = 0;
    assign rom[13'h1fb7] = 0;
    assign rom[13'h1fb8] = 0;
    assign rom[13'h1fb9] = 0;
    assign rom[13'h1fba] = 0;
    assign rom[13'h1fbb] = 0;
    assign rom[13'h1fbc] = 0;
    assign rom[13'h1fbd] = 0;
    assign rom[13'h1fbe] = 0;
    assign rom[13'h1fbf] = 0;
    assign rom[13'h1fc0] = 1;
    assign rom[13'h1fc1] = 1;
    assign rom[13'h1fc2] = 1;
    assign rom[13'h1fc3] = 1;
    assign rom[13'h1fc4] = 1;
    assign rom[13'h1fc5] = 1;
    assign rom[13'h1fc6] = 1;
    assign rom[13'h1fc7] = 1;
    assign rom[13'h1fc8] = 1;
    assign rom[13'h1fc9] = 1;
    assign rom[13'h1fca] = 1;
    assign rom[13'h1fcb] = 1;
    assign rom[13'h1fcc] = 1;
    assign rom[13'h1fcd] = 1;
    assign rom[13'h1fce] = 1;
    assign rom[13'h1fcf] = 1;
    assign rom[13'h1fd0] = 1;
    assign rom[13'h1fd1] = 1;
    assign rom[13'h1fd2] = 1;
    assign rom[13'h1fd3] = 1;
    assign rom[13'h1fd4] = 1;
    assign rom[13'h1fd5] = 1;
    assign rom[13'h1fd6] = 1;
    assign rom[13'h1fd7] = 1;
    assign rom[13'h1fd8] = 1;
    assign rom[13'h1fd9] = 1;
    assign rom[13'h1fda] = 1;
    assign rom[13'h1fdb] = 1;
    assign rom[13'h1fdc] = 1;
    assign rom[13'h1fdd] = 1;
    assign rom[13'h1fde] = 1;
    assign rom[13'h1fdf] = 1;
    assign rom[13'h1fe0] = 1;
    assign rom[13'h1fe1] = 1;
    assign rom[13'h1fe2] = 1;
    assign rom[13'h1fe3] = 1;
    assign rom[13'h1fe4] = 1;
    assign rom[13'h1fe5] = 1;
    assign rom[13'h1fe6] = 1;
    assign rom[13'h1fe7] = 1;
    assign rom[13'h1fe8] = 1;
    assign rom[13'h1fe9] = 1;
    assign rom[13'h1fea] = 1;
    assign rom[13'h1feb] = 1;
    assign rom[13'h1fec] = 1;
    assign rom[13'h1fed] = 1;
    assign rom[13'h1fee] = 1;
    assign rom[13'h1fef] = 1;
    assign rom[13'h1ff0] = 1;
    assign rom[13'h1ff1] = 1;
    assign rom[13'h1ff2] = 1;
    assign rom[13'h1ff3] = 1;
    assign rom[13'h1ff4] = 1;
    assign rom[13'h1ff5] = 1;
    assign rom[13'h1ff6] = 1;
    assign rom[13'h1ff7] = 1;
    assign rom[13'h1ff8] = 1;
    assign rom[13'h1ff9] = 1;
    assign rom[13'h1ffa] = 1;
    assign rom[13'h1ffb] = 1;
    assign rom[13'h1ffc] = 1;
    assign rom[13'h1ffd] = 1;
    assign rom[13'h1ffe] = 1;
    assign rom[13'h1fff] = 1;
endmodule
